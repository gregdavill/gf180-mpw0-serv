// This is the unpowered netlist.
module serv_1 (io_in,
    io_oeb,
    io_out);
 input [4:0] io_in;
 output [4:0] io_oeb;
 output [4:0] io_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire \u_arbiter.i_wb_cpu_ack ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[10] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[11] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[12] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[13] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[14] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[15] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[16] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[17] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[18] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[19] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[20] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[21] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[22] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[23] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[24] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[25] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[26] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[27] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[28] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[29] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[2] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[30] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[31] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[3] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[4] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[5] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[6] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[7] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[8] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[9] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[0] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[10] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[11] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[12] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[13] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[14] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[15] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[16] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[17] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[18] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[19] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[1] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[20] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[21] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[22] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[23] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[24] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[25] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[26] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[27] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[28] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[29] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[2] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[30] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[31] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[3] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[4] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[5] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[6] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[7] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[8] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[9] ;
 wire \u_arbiter.i_wb_cpu_dbus_sel[0] ;
 wire \u_arbiter.i_wb_cpu_dbus_sel[1] ;
 wire \u_arbiter.i_wb_cpu_dbus_sel[2] ;
 wire \u_arbiter.i_wb_cpu_dbus_sel[3] ;
 wire \u_arbiter.i_wb_cpu_dbus_we ;
 wire \u_arbiter.i_wb_cpu_ibus_adr[0] ;
 wire \u_arbiter.i_wb_cpu_ibus_adr[1] ;
 wire \u_arbiter.i_wb_cpu_rdt[0] ;
 wire \u_arbiter.i_wb_cpu_rdt[10] ;
 wire \u_arbiter.i_wb_cpu_rdt[11] ;
 wire \u_arbiter.i_wb_cpu_rdt[12] ;
 wire \u_arbiter.i_wb_cpu_rdt[13] ;
 wire \u_arbiter.i_wb_cpu_rdt[14] ;
 wire \u_arbiter.i_wb_cpu_rdt[15] ;
 wire \u_arbiter.i_wb_cpu_rdt[16] ;
 wire \u_arbiter.i_wb_cpu_rdt[17] ;
 wire \u_arbiter.i_wb_cpu_rdt[18] ;
 wire \u_arbiter.i_wb_cpu_rdt[19] ;
 wire \u_arbiter.i_wb_cpu_rdt[1] ;
 wire \u_arbiter.i_wb_cpu_rdt[20] ;
 wire \u_arbiter.i_wb_cpu_rdt[21] ;
 wire \u_arbiter.i_wb_cpu_rdt[22] ;
 wire \u_arbiter.i_wb_cpu_rdt[23] ;
 wire \u_arbiter.i_wb_cpu_rdt[24] ;
 wire \u_arbiter.i_wb_cpu_rdt[25] ;
 wire \u_arbiter.i_wb_cpu_rdt[26] ;
 wire \u_arbiter.i_wb_cpu_rdt[27] ;
 wire \u_arbiter.i_wb_cpu_rdt[28] ;
 wire \u_arbiter.i_wb_cpu_rdt[29] ;
 wire \u_arbiter.i_wb_cpu_rdt[2] ;
 wire \u_arbiter.i_wb_cpu_rdt[30] ;
 wire \u_arbiter.i_wb_cpu_rdt[31] ;
 wire \u_arbiter.i_wb_cpu_rdt[3] ;
 wire \u_arbiter.i_wb_cpu_rdt[4] ;
 wire \u_arbiter.i_wb_cpu_rdt[5] ;
 wire \u_arbiter.i_wb_cpu_rdt[6] ;
 wire \u_arbiter.i_wb_cpu_rdt[7] ;
 wire \u_arbiter.i_wb_cpu_rdt[8] ;
 wire \u_arbiter.i_wb_cpu_rdt[9] ;
 wire \u_arbiter.o_wb_cpu_adr[0] ;
 wire \u_arbiter.o_wb_cpu_adr[10] ;
 wire \u_arbiter.o_wb_cpu_adr[11] ;
 wire \u_arbiter.o_wb_cpu_adr[12] ;
 wire \u_arbiter.o_wb_cpu_adr[13] ;
 wire \u_arbiter.o_wb_cpu_adr[14] ;
 wire \u_arbiter.o_wb_cpu_adr[15] ;
 wire \u_arbiter.o_wb_cpu_adr[16] ;
 wire \u_arbiter.o_wb_cpu_adr[17] ;
 wire \u_arbiter.o_wb_cpu_adr[18] ;
 wire \u_arbiter.o_wb_cpu_adr[19] ;
 wire \u_arbiter.o_wb_cpu_adr[1] ;
 wire \u_arbiter.o_wb_cpu_adr[20] ;
 wire \u_arbiter.o_wb_cpu_adr[21] ;
 wire \u_arbiter.o_wb_cpu_adr[22] ;
 wire \u_arbiter.o_wb_cpu_adr[23] ;
 wire \u_arbiter.o_wb_cpu_adr[24] ;
 wire \u_arbiter.o_wb_cpu_adr[25] ;
 wire \u_arbiter.o_wb_cpu_adr[26] ;
 wire \u_arbiter.o_wb_cpu_adr[27] ;
 wire \u_arbiter.o_wb_cpu_adr[28] ;
 wire \u_arbiter.o_wb_cpu_adr[29] ;
 wire \u_arbiter.o_wb_cpu_adr[2] ;
 wire \u_arbiter.o_wb_cpu_adr[30] ;
 wire \u_arbiter.o_wb_cpu_adr[31] ;
 wire \u_arbiter.o_wb_cpu_adr[3] ;
 wire \u_arbiter.o_wb_cpu_adr[4] ;
 wire \u_arbiter.o_wb_cpu_adr[5] ;
 wire \u_arbiter.o_wb_cpu_adr[6] ;
 wire \u_arbiter.o_wb_cpu_adr[7] ;
 wire \u_arbiter.o_wb_cpu_adr[8] ;
 wire \u_arbiter.o_wb_cpu_adr[9] ;
 wire \u_arbiter.o_wb_cpu_cyc ;
 wire \u_arbiter.o_wb_cpu_we ;
 wire \u_cpu.cpu.alu.add_cy_r ;
 wire \u_cpu.cpu.alu.cmp_r ;
 wire \u_cpu.cpu.alu.i_rs1 ;
 wire \u_cpu.cpu.bne_or_bge ;
 wire \u_cpu.cpu.branch_op ;
 wire \u_cpu.cpu.bufreg.c_r ;
 wire \u_cpu.cpu.bufreg.i_sh_signed ;
 wire \u_cpu.cpu.bufreg.lsb[0] ;
 wire \u_cpu.cpu.bufreg.lsb[1] ;
 wire \u_cpu.cpu.bufreg2.i_cnt_done ;
 wire \u_cpu.cpu.csr_d_sel ;
 wire \u_cpu.cpu.csr_imm ;
 wire \u_cpu.cpu.ctrl.i_iscomp ;
 wire \u_cpu.cpu.ctrl.i_jump ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[10] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[11] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[12] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[13] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[14] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[15] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[16] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[17] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[18] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[19] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[20] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[21] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[22] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[23] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[24] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[25] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[26] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[27] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[28] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[29] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[2] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[30] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[31] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[3] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[4] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[5] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[6] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[7] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[8] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[9] ;
 wire \u_cpu.cpu.ctrl.pc_plus_4_cy_r ;
 wire \u_cpu.cpu.ctrl.pc_plus_offset_cy_r ;
 wire \u_cpu.cpu.decode.co_ebreak ;
 wire \u_cpu.cpu.decode.co_mem_word ;
 wire \u_cpu.cpu.decode.op21 ;
 wire \u_cpu.cpu.decode.op22 ;
 wire \u_cpu.cpu.decode.op26 ;
 wire \u_cpu.cpu.decode.opcode[0] ;
 wire \u_cpu.cpu.decode.opcode[1] ;
 wire \u_cpu.cpu.decode.opcode[2] ;
 wire \u_cpu.cpu.genblk1.align.ctrl_misal ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[10] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[11] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[2] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[3] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ;
 wire \u_cpu.cpu.genblk3.csr.i_mtip ;
 wire \u_cpu.cpu.genblk3.csr.mcause31 ;
 wire \u_cpu.cpu.genblk3.csr.mcause3_0[0] ;
 wire \u_cpu.cpu.genblk3.csr.mcause3_0[1] ;
 wire \u_cpu.cpu.genblk3.csr.mcause3_0[2] ;
 wire \u_cpu.cpu.genblk3.csr.mcause3_0[3] ;
 wire \u_cpu.cpu.genblk3.csr.mie_mtie ;
 wire \u_cpu.cpu.genblk3.csr.mstatus_mie ;
 wire \u_cpu.cpu.genblk3.csr.mstatus_mpie ;
 wire \u_cpu.cpu.genblk3.csr.o_new_irq ;
 wire \u_cpu.cpu.genblk3.csr.timer_irq_r ;
 wire \u_cpu.cpu.immdec.imm11_7[0] ;
 wire \u_cpu.cpu.immdec.imm11_7[1] ;
 wire \u_cpu.cpu.immdec.imm11_7[2] ;
 wire \u_cpu.cpu.immdec.imm11_7[3] ;
 wire \u_cpu.cpu.immdec.imm11_7[4] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[0] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[1] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[2] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[3] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[5] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[6] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[7] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[8] ;
 wire \u_cpu.cpu.immdec.imm24_20[0] ;
 wire \u_cpu.cpu.immdec.imm24_20[1] ;
 wire \u_cpu.cpu.immdec.imm24_20[2] ;
 wire \u_cpu.cpu.immdec.imm24_20[3] ;
 wire \u_cpu.cpu.immdec.imm24_20[4] ;
 wire \u_cpu.cpu.immdec.imm30_25[0] ;
 wire \u_cpu.cpu.immdec.imm30_25[1] ;
 wire \u_cpu.cpu.immdec.imm30_25[2] ;
 wire \u_cpu.cpu.immdec.imm30_25[3] ;
 wire \u_cpu.cpu.immdec.imm30_25[4] ;
 wire \u_cpu.cpu.immdec.imm30_25[5] ;
 wire \u_cpu.cpu.immdec.imm31 ;
 wire \u_cpu.cpu.immdec.imm7 ;
 wire \u_cpu.cpu.mem_bytecnt[0] ;
 wire \u_cpu.cpu.mem_bytecnt[1] ;
 wire \u_cpu.cpu.mem_if.signbit ;
 wire \u_cpu.cpu.o_wdata0 ;
 wire \u_cpu.cpu.o_wdata1 ;
 wire \u_cpu.cpu.o_wen0 ;
 wire \u_cpu.cpu.o_wen1 ;
 wire \u_cpu.cpu.state.genblk1.misalign_trap_sync_r ;
 wire \u_cpu.cpu.state.ibus_cyc ;
 wire \u_cpu.cpu.state.init_done ;
 wire \u_cpu.cpu.state.o_cnt[2] ;
 wire \u_cpu.cpu.state.o_cnt_r[0] ;
 wire \u_cpu.cpu.state.o_cnt_r[1] ;
 wire \u_cpu.cpu.state.o_cnt_r[2] ;
 wire \u_cpu.cpu.state.o_cnt_r[3] ;
 wire \u_cpu.cpu.state.stage_two_req ;
 wire \u_cpu.raddr[0] ;
 wire \u_cpu.raddr[1] ;
 wire \u_cpu.rf_ram.memory[0][0] ;
 wire \u_cpu.rf_ram.memory[0][1] ;
 wire \u_cpu.rf_ram.memory[0][2] ;
 wire \u_cpu.rf_ram.memory[0][3] ;
 wire \u_cpu.rf_ram.memory[0][4] ;
 wire \u_cpu.rf_ram.memory[0][5] ;
 wire \u_cpu.rf_ram.memory[0][6] ;
 wire \u_cpu.rf_ram.memory[0][7] ;
 wire \u_cpu.rf_ram.memory[100][0] ;
 wire \u_cpu.rf_ram.memory[100][1] ;
 wire \u_cpu.rf_ram.memory[100][2] ;
 wire \u_cpu.rf_ram.memory[100][3] ;
 wire \u_cpu.rf_ram.memory[100][4] ;
 wire \u_cpu.rf_ram.memory[100][5] ;
 wire \u_cpu.rf_ram.memory[100][6] ;
 wire \u_cpu.rf_ram.memory[100][7] ;
 wire \u_cpu.rf_ram.memory[101][0] ;
 wire \u_cpu.rf_ram.memory[101][1] ;
 wire \u_cpu.rf_ram.memory[101][2] ;
 wire \u_cpu.rf_ram.memory[101][3] ;
 wire \u_cpu.rf_ram.memory[101][4] ;
 wire \u_cpu.rf_ram.memory[101][5] ;
 wire \u_cpu.rf_ram.memory[101][6] ;
 wire \u_cpu.rf_ram.memory[101][7] ;
 wire \u_cpu.rf_ram.memory[102][0] ;
 wire \u_cpu.rf_ram.memory[102][1] ;
 wire \u_cpu.rf_ram.memory[102][2] ;
 wire \u_cpu.rf_ram.memory[102][3] ;
 wire \u_cpu.rf_ram.memory[102][4] ;
 wire \u_cpu.rf_ram.memory[102][5] ;
 wire \u_cpu.rf_ram.memory[102][6] ;
 wire \u_cpu.rf_ram.memory[102][7] ;
 wire \u_cpu.rf_ram.memory[103][0] ;
 wire \u_cpu.rf_ram.memory[103][1] ;
 wire \u_cpu.rf_ram.memory[103][2] ;
 wire \u_cpu.rf_ram.memory[103][3] ;
 wire \u_cpu.rf_ram.memory[103][4] ;
 wire \u_cpu.rf_ram.memory[103][5] ;
 wire \u_cpu.rf_ram.memory[103][6] ;
 wire \u_cpu.rf_ram.memory[103][7] ;
 wire \u_cpu.rf_ram.memory[104][0] ;
 wire \u_cpu.rf_ram.memory[104][1] ;
 wire \u_cpu.rf_ram.memory[104][2] ;
 wire \u_cpu.rf_ram.memory[104][3] ;
 wire \u_cpu.rf_ram.memory[104][4] ;
 wire \u_cpu.rf_ram.memory[104][5] ;
 wire \u_cpu.rf_ram.memory[104][6] ;
 wire \u_cpu.rf_ram.memory[104][7] ;
 wire \u_cpu.rf_ram.memory[105][0] ;
 wire \u_cpu.rf_ram.memory[105][1] ;
 wire \u_cpu.rf_ram.memory[105][2] ;
 wire \u_cpu.rf_ram.memory[105][3] ;
 wire \u_cpu.rf_ram.memory[105][4] ;
 wire \u_cpu.rf_ram.memory[105][5] ;
 wire \u_cpu.rf_ram.memory[105][6] ;
 wire \u_cpu.rf_ram.memory[105][7] ;
 wire \u_cpu.rf_ram.memory[106][0] ;
 wire \u_cpu.rf_ram.memory[106][1] ;
 wire \u_cpu.rf_ram.memory[106][2] ;
 wire \u_cpu.rf_ram.memory[106][3] ;
 wire \u_cpu.rf_ram.memory[106][4] ;
 wire \u_cpu.rf_ram.memory[106][5] ;
 wire \u_cpu.rf_ram.memory[106][6] ;
 wire \u_cpu.rf_ram.memory[106][7] ;
 wire \u_cpu.rf_ram.memory[107][0] ;
 wire \u_cpu.rf_ram.memory[107][1] ;
 wire \u_cpu.rf_ram.memory[107][2] ;
 wire \u_cpu.rf_ram.memory[107][3] ;
 wire \u_cpu.rf_ram.memory[107][4] ;
 wire \u_cpu.rf_ram.memory[107][5] ;
 wire \u_cpu.rf_ram.memory[107][6] ;
 wire \u_cpu.rf_ram.memory[107][7] ;
 wire \u_cpu.rf_ram.memory[108][0] ;
 wire \u_cpu.rf_ram.memory[108][1] ;
 wire \u_cpu.rf_ram.memory[108][2] ;
 wire \u_cpu.rf_ram.memory[108][3] ;
 wire \u_cpu.rf_ram.memory[108][4] ;
 wire \u_cpu.rf_ram.memory[108][5] ;
 wire \u_cpu.rf_ram.memory[108][6] ;
 wire \u_cpu.rf_ram.memory[108][7] ;
 wire \u_cpu.rf_ram.memory[109][0] ;
 wire \u_cpu.rf_ram.memory[109][1] ;
 wire \u_cpu.rf_ram.memory[109][2] ;
 wire \u_cpu.rf_ram.memory[109][3] ;
 wire \u_cpu.rf_ram.memory[109][4] ;
 wire \u_cpu.rf_ram.memory[109][5] ;
 wire \u_cpu.rf_ram.memory[109][6] ;
 wire \u_cpu.rf_ram.memory[109][7] ;
 wire \u_cpu.rf_ram.memory[10][0] ;
 wire \u_cpu.rf_ram.memory[10][1] ;
 wire \u_cpu.rf_ram.memory[10][2] ;
 wire \u_cpu.rf_ram.memory[10][3] ;
 wire \u_cpu.rf_ram.memory[10][4] ;
 wire \u_cpu.rf_ram.memory[10][5] ;
 wire \u_cpu.rf_ram.memory[10][6] ;
 wire \u_cpu.rf_ram.memory[10][7] ;
 wire \u_cpu.rf_ram.memory[110][0] ;
 wire \u_cpu.rf_ram.memory[110][1] ;
 wire \u_cpu.rf_ram.memory[110][2] ;
 wire \u_cpu.rf_ram.memory[110][3] ;
 wire \u_cpu.rf_ram.memory[110][4] ;
 wire \u_cpu.rf_ram.memory[110][5] ;
 wire \u_cpu.rf_ram.memory[110][6] ;
 wire \u_cpu.rf_ram.memory[110][7] ;
 wire \u_cpu.rf_ram.memory[111][0] ;
 wire \u_cpu.rf_ram.memory[111][1] ;
 wire \u_cpu.rf_ram.memory[111][2] ;
 wire \u_cpu.rf_ram.memory[111][3] ;
 wire \u_cpu.rf_ram.memory[111][4] ;
 wire \u_cpu.rf_ram.memory[111][5] ;
 wire \u_cpu.rf_ram.memory[111][6] ;
 wire \u_cpu.rf_ram.memory[111][7] ;
 wire \u_cpu.rf_ram.memory[112][0] ;
 wire \u_cpu.rf_ram.memory[112][1] ;
 wire \u_cpu.rf_ram.memory[112][2] ;
 wire \u_cpu.rf_ram.memory[112][3] ;
 wire \u_cpu.rf_ram.memory[112][4] ;
 wire \u_cpu.rf_ram.memory[112][5] ;
 wire \u_cpu.rf_ram.memory[112][6] ;
 wire \u_cpu.rf_ram.memory[112][7] ;
 wire \u_cpu.rf_ram.memory[113][0] ;
 wire \u_cpu.rf_ram.memory[113][1] ;
 wire \u_cpu.rf_ram.memory[113][2] ;
 wire \u_cpu.rf_ram.memory[113][3] ;
 wire \u_cpu.rf_ram.memory[113][4] ;
 wire \u_cpu.rf_ram.memory[113][5] ;
 wire \u_cpu.rf_ram.memory[113][6] ;
 wire \u_cpu.rf_ram.memory[113][7] ;
 wire \u_cpu.rf_ram.memory[114][0] ;
 wire \u_cpu.rf_ram.memory[114][1] ;
 wire \u_cpu.rf_ram.memory[114][2] ;
 wire \u_cpu.rf_ram.memory[114][3] ;
 wire \u_cpu.rf_ram.memory[114][4] ;
 wire \u_cpu.rf_ram.memory[114][5] ;
 wire \u_cpu.rf_ram.memory[114][6] ;
 wire \u_cpu.rf_ram.memory[114][7] ;
 wire \u_cpu.rf_ram.memory[115][0] ;
 wire \u_cpu.rf_ram.memory[115][1] ;
 wire \u_cpu.rf_ram.memory[115][2] ;
 wire \u_cpu.rf_ram.memory[115][3] ;
 wire \u_cpu.rf_ram.memory[115][4] ;
 wire \u_cpu.rf_ram.memory[115][5] ;
 wire \u_cpu.rf_ram.memory[115][6] ;
 wire \u_cpu.rf_ram.memory[115][7] ;
 wire \u_cpu.rf_ram.memory[116][0] ;
 wire \u_cpu.rf_ram.memory[116][1] ;
 wire \u_cpu.rf_ram.memory[116][2] ;
 wire \u_cpu.rf_ram.memory[116][3] ;
 wire \u_cpu.rf_ram.memory[116][4] ;
 wire \u_cpu.rf_ram.memory[116][5] ;
 wire \u_cpu.rf_ram.memory[116][6] ;
 wire \u_cpu.rf_ram.memory[116][7] ;
 wire \u_cpu.rf_ram.memory[117][0] ;
 wire \u_cpu.rf_ram.memory[117][1] ;
 wire \u_cpu.rf_ram.memory[117][2] ;
 wire \u_cpu.rf_ram.memory[117][3] ;
 wire \u_cpu.rf_ram.memory[117][4] ;
 wire \u_cpu.rf_ram.memory[117][5] ;
 wire \u_cpu.rf_ram.memory[117][6] ;
 wire \u_cpu.rf_ram.memory[117][7] ;
 wire \u_cpu.rf_ram.memory[118][0] ;
 wire \u_cpu.rf_ram.memory[118][1] ;
 wire \u_cpu.rf_ram.memory[118][2] ;
 wire \u_cpu.rf_ram.memory[118][3] ;
 wire \u_cpu.rf_ram.memory[118][4] ;
 wire \u_cpu.rf_ram.memory[118][5] ;
 wire \u_cpu.rf_ram.memory[118][6] ;
 wire \u_cpu.rf_ram.memory[118][7] ;
 wire \u_cpu.rf_ram.memory[119][0] ;
 wire \u_cpu.rf_ram.memory[119][1] ;
 wire \u_cpu.rf_ram.memory[119][2] ;
 wire \u_cpu.rf_ram.memory[119][3] ;
 wire \u_cpu.rf_ram.memory[119][4] ;
 wire \u_cpu.rf_ram.memory[119][5] ;
 wire \u_cpu.rf_ram.memory[119][6] ;
 wire \u_cpu.rf_ram.memory[119][7] ;
 wire \u_cpu.rf_ram.memory[11][0] ;
 wire \u_cpu.rf_ram.memory[11][1] ;
 wire \u_cpu.rf_ram.memory[11][2] ;
 wire \u_cpu.rf_ram.memory[11][3] ;
 wire \u_cpu.rf_ram.memory[11][4] ;
 wire \u_cpu.rf_ram.memory[11][5] ;
 wire \u_cpu.rf_ram.memory[11][6] ;
 wire \u_cpu.rf_ram.memory[11][7] ;
 wire \u_cpu.rf_ram.memory[120][0] ;
 wire \u_cpu.rf_ram.memory[120][1] ;
 wire \u_cpu.rf_ram.memory[120][2] ;
 wire \u_cpu.rf_ram.memory[120][3] ;
 wire \u_cpu.rf_ram.memory[120][4] ;
 wire \u_cpu.rf_ram.memory[120][5] ;
 wire \u_cpu.rf_ram.memory[120][6] ;
 wire \u_cpu.rf_ram.memory[120][7] ;
 wire \u_cpu.rf_ram.memory[121][0] ;
 wire \u_cpu.rf_ram.memory[121][1] ;
 wire \u_cpu.rf_ram.memory[121][2] ;
 wire \u_cpu.rf_ram.memory[121][3] ;
 wire \u_cpu.rf_ram.memory[121][4] ;
 wire \u_cpu.rf_ram.memory[121][5] ;
 wire \u_cpu.rf_ram.memory[121][6] ;
 wire \u_cpu.rf_ram.memory[121][7] ;
 wire \u_cpu.rf_ram.memory[122][0] ;
 wire \u_cpu.rf_ram.memory[122][1] ;
 wire \u_cpu.rf_ram.memory[122][2] ;
 wire \u_cpu.rf_ram.memory[122][3] ;
 wire \u_cpu.rf_ram.memory[122][4] ;
 wire \u_cpu.rf_ram.memory[122][5] ;
 wire \u_cpu.rf_ram.memory[122][6] ;
 wire \u_cpu.rf_ram.memory[122][7] ;
 wire \u_cpu.rf_ram.memory[123][0] ;
 wire \u_cpu.rf_ram.memory[123][1] ;
 wire \u_cpu.rf_ram.memory[123][2] ;
 wire \u_cpu.rf_ram.memory[123][3] ;
 wire \u_cpu.rf_ram.memory[123][4] ;
 wire \u_cpu.rf_ram.memory[123][5] ;
 wire \u_cpu.rf_ram.memory[123][6] ;
 wire \u_cpu.rf_ram.memory[123][7] ;
 wire \u_cpu.rf_ram.memory[124][0] ;
 wire \u_cpu.rf_ram.memory[124][1] ;
 wire \u_cpu.rf_ram.memory[124][2] ;
 wire \u_cpu.rf_ram.memory[124][3] ;
 wire \u_cpu.rf_ram.memory[124][4] ;
 wire \u_cpu.rf_ram.memory[124][5] ;
 wire \u_cpu.rf_ram.memory[124][6] ;
 wire \u_cpu.rf_ram.memory[124][7] ;
 wire \u_cpu.rf_ram.memory[125][0] ;
 wire \u_cpu.rf_ram.memory[125][1] ;
 wire \u_cpu.rf_ram.memory[125][2] ;
 wire \u_cpu.rf_ram.memory[125][3] ;
 wire \u_cpu.rf_ram.memory[125][4] ;
 wire \u_cpu.rf_ram.memory[125][5] ;
 wire \u_cpu.rf_ram.memory[125][6] ;
 wire \u_cpu.rf_ram.memory[125][7] ;
 wire \u_cpu.rf_ram.memory[126][0] ;
 wire \u_cpu.rf_ram.memory[126][1] ;
 wire \u_cpu.rf_ram.memory[126][2] ;
 wire \u_cpu.rf_ram.memory[126][3] ;
 wire \u_cpu.rf_ram.memory[126][4] ;
 wire \u_cpu.rf_ram.memory[126][5] ;
 wire \u_cpu.rf_ram.memory[126][6] ;
 wire \u_cpu.rf_ram.memory[126][7] ;
 wire \u_cpu.rf_ram.memory[127][0] ;
 wire \u_cpu.rf_ram.memory[127][1] ;
 wire \u_cpu.rf_ram.memory[127][2] ;
 wire \u_cpu.rf_ram.memory[127][3] ;
 wire \u_cpu.rf_ram.memory[127][4] ;
 wire \u_cpu.rf_ram.memory[127][5] ;
 wire \u_cpu.rf_ram.memory[127][6] ;
 wire \u_cpu.rf_ram.memory[127][7] ;
 wire \u_cpu.rf_ram.memory[128][0] ;
 wire \u_cpu.rf_ram.memory[128][1] ;
 wire \u_cpu.rf_ram.memory[128][2] ;
 wire \u_cpu.rf_ram.memory[128][3] ;
 wire \u_cpu.rf_ram.memory[128][4] ;
 wire \u_cpu.rf_ram.memory[128][5] ;
 wire \u_cpu.rf_ram.memory[128][6] ;
 wire \u_cpu.rf_ram.memory[128][7] ;
 wire \u_cpu.rf_ram.memory[129][0] ;
 wire \u_cpu.rf_ram.memory[129][1] ;
 wire \u_cpu.rf_ram.memory[129][2] ;
 wire \u_cpu.rf_ram.memory[129][3] ;
 wire \u_cpu.rf_ram.memory[129][4] ;
 wire \u_cpu.rf_ram.memory[129][5] ;
 wire \u_cpu.rf_ram.memory[129][6] ;
 wire \u_cpu.rf_ram.memory[129][7] ;
 wire \u_cpu.rf_ram.memory[12][0] ;
 wire \u_cpu.rf_ram.memory[12][1] ;
 wire \u_cpu.rf_ram.memory[12][2] ;
 wire \u_cpu.rf_ram.memory[12][3] ;
 wire \u_cpu.rf_ram.memory[12][4] ;
 wire \u_cpu.rf_ram.memory[12][5] ;
 wire \u_cpu.rf_ram.memory[12][6] ;
 wire \u_cpu.rf_ram.memory[12][7] ;
 wire \u_cpu.rf_ram.memory[130][0] ;
 wire \u_cpu.rf_ram.memory[130][1] ;
 wire \u_cpu.rf_ram.memory[130][2] ;
 wire \u_cpu.rf_ram.memory[130][3] ;
 wire \u_cpu.rf_ram.memory[130][4] ;
 wire \u_cpu.rf_ram.memory[130][5] ;
 wire \u_cpu.rf_ram.memory[130][6] ;
 wire \u_cpu.rf_ram.memory[130][7] ;
 wire \u_cpu.rf_ram.memory[131][0] ;
 wire \u_cpu.rf_ram.memory[131][1] ;
 wire \u_cpu.rf_ram.memory[131][2] ;
 wire \u_cpu.rf_ram.memory[131][3] ;
 wire \u_cpu.rf_ram.memory[131][4] ;
 wire \u_cpu.rf_ram.memory[131][5] ;
 wire \u_cpu.rf_ram.memory[131][6] ;
 wire \u_cpu.rf_ram.memory[131][7] ;
 wire \u_cpu.rf_ram.memory[132][0] ;
 wire \u_cpu.rf_ram.memory[132][1] ;
 wire \u_cpu.rf_ram.memory[132][2] ;
 wire \u_cpu.rf_ram.memory[132][3] ;
 wire \u_cpu.rf_ram.memory[132][4] ;
 wire \u_cpu.rf_ram.memory[132][5] ;
 wire \u_cpu.rf_ram.memory[132][6] ;
 wire \u_cpu.rf_ram.memory[132][7] ;
 wire \u_cpu.rf_ram.memory[133][0] ;
 wire \u_cpu.rf_ram.memory[133][1] ;
 wire \u_cpu.rf_ram.memory[133][2] ;
 wire \u_cpu.rf_ram.memory[133][3] ;
 wire \u_cpu.rf_ram.memory[133][4] ;
 wire \u_cpu.rf_ram.memory[133][5] ;
 wire \u_cpu.rf_ram.memory[133][6] ;
 wire \u_cpu.rf_ram.memory[133][7] ;
 wire \u_cpu.rf_ram.memory[134][0] ;
 wire \u_cpu.rf_ram.memory[134][1] ;
 wire \u_cpu.rf_ram.memory[134][2] ;
 wire \u_cpu.rf_ram.memory[134][3] ;
 wire \u_cpu.rf_ram.memory[134][4] ;
 wire \u_cpu.rf_ram.memory[134][5] ;
 wire \u_cpu.rf_ram.memory[134][6] ;
 wire \u_cpu.rf_ram.memory[134][7] ;
 wire \u_cpu.rf_ram.memory[135][0] ;
 wire \u_cpu.rf_ram.memory[135][1] ;
 wire \u_cpu.rf_ram.memory[135][2] ;
 wire \u_cpu.rf_ram.memory[135][3] ;
 wire \u_cpu.rf_ram.memory[135][4] ;
 wire \u_cpu.rf_ram.memory[135][5] ;
 wire \u_cpu.rf_ram.memory[135][6] ;
 wire \u_cpu.rf_ram.memory[135][7] ;
 wire \u_cpu.rf_ram.memory[136][0] ;
 wire \u_cpu.rf_ram.memory[136][1] ;
 wire \u_cpu.rf_ram.memory[136][2] ;
 wire \u_cpu.rf_ram.memory[136][3] ;
 wire \u_cpu.rf_ram.memory[136][4] ;
 wire \u_cpu.rf_ram.memory[136][5] ;
 wire \u_cpu.rf_ram.memory[136][6] ;
 wire \u_cpu.rf_ram.memory[136][7] ;
 wire \u_cpu.rf_ram.memory[137][0] ;
 wire \u_cpu.rf_ram.memory[137][1] ;
 wire \u_cpu.rf_ram.memory[137][2] ;
 wire \u_cpu.rf_ram.memory[137][3] ;
 wire \u_cpu.rf_ram.memory[137][4] ;
 wire \u_cpu.rf_ram.memory[137][5] ;
 wire \u_cpu.rf_ram.memory[137][6] ;
 wire \u_cpu.rf_ram.memory[137][7] ;
 wire \u_cpu.rf_ram.memory[138][0] ;
 wire \u_cpu.rf_ram.memory[138][1] ;
 wire \u_cpu.rf_ram.memory[138][2] ;
 wire \u_cpu.rf_ram.memory[138][3] ;
 wire \u_cpu.rf_ram.memory[138][4] ;
 wire \u_cpu.rf_ram.memory[138][5] ;
 wire \u_cpu.rf_ram.memory[138][6] ;
 wire \u_cpu.rf_ram.memory[138][7] ;
 wire \u_cpu.rf_ram.memory[139][0] ;
 wire \u_cpu.rf_ram.memory[139][1] ;
 wire \u_cpu.rf_ram.memory[139][2] ;
 wire \u_cpu.rf_ram.memory[139][3] ;
 wire \u_cpu.rf_ram.memory[139][4] ;
 wire \u_cpu.rf_ram.memory[139][5] ;
 wire \u_cpu.rf_ram.memory[139][6] ;
 wire \u_cpu.rf_ram.memory[139][7] ;
 wire \u_cpu.rf_ram.memory[13][0] ;
 wire \u_cpu.rf_ram.memory[13][1] ;
 wire \u_cpu.rf_ram.memory[13][2] ;
 wire \u_cpu.rf_ram.memory[13][3] ;
 wire \u_cpu.rf_ram.memory[13][4] ;
 wire \u_cpu.rf_ram.memory[13][5] ;
 wire \u_cpu.rf_ram.memory[13][6] ;
 wire \u_cpu.rf_ram.memory[13][7] ;
 wire \u_cpu.rf_ram.memory[140][0] ;
 wire \u_cpu.rf_ram.memory[140][1] ;
 wire \u_cpu.rf_ram.memory[140][2] ;
 wire \u_cpu.rf_ram.memory[140][3] ;
 wire \u_cpu.rf_ram.memory[140][4] ;
 wire \u_cpu.rf_ram.memory[140][5] ;
 wire \u_cpu.rf_ram.memory[140][6] ;
 wire \u_cpu.rf_ram.memory[140][7] ;
 wire \u_cpu.rf_ram.memory[141][0] ;
 wire \u_cpu.rf_ram.memory[141][1] ;
 wire \u_cpu.rf_ram.memory[141][2] ;
 wire \u_cpu.rf_ram.memory[141][3] ;
 wire \u_cpu.rf_ram.memory[141][4] ;
 wire \u_cpu.rf_ram.memory[141][5] ;
 wire \u_cpu.rf_ram.memory[141][6] ;
 wire \u_cpu.rf_ram.memory[141][7] ;
 wire \u_cpu.rf_ram.memory[142][0] ;
 wire \u_cpu.rf_ram.memory[142][1] ;
 wire \u_cpu.rf_ram.memory[142][2] ;
 wire \u_cpu.rf_ram.memory[142][3] ;
 wire \u_cpu.rf_ram.memory[142][4] ;
 wire \u_cpu.rf_ram.memory[142][5] ;
 wire \u_cpu.rf_ram.memory[142][6] ;
 wire \u_cpu.rf_ram.memory[142][7] ;
 wire \u_cpu.rf_ram.memory[143][0] ;
 wire \u_cpu.rf_ram.memory[143][1] ;
 wire \u_cpu.rf_ram.memory[143][2] ;
 wire \u_cpu.rf_ram.memory[143][3] ;
 wire \u_cpu.rf_ram.memory[143][4] ;
 wire \u_cpu.rf_ram.memory[143][5] ;
 wire \u_cpu.rf_ram.memory[143][6] ;
 wire \u_cpu.rf_ram.memory[143][7] ;
 wire \u_cpu.rf_ram.memory[14][0] ;
 wire \u_cpu.rf_ram.memory[14][1] ;
 wire \u_cpu.rf_ram.memory[14][2] ;
 wire \u_cpu.rf_ram.memory[14][3] ;
 wire \u_cpu.rf_ram.memory[14][4] ;
 wire \u_cpu.rf_ram.memory[14][5] ;
 wire \u_cpu.rf_ram.memory[14][6] ;
 wire \u_cpu.rf_ram.memory[14][7] ;
 wire \u_cpu.rf_ram.memory[15][0] ;
 wire \u_cpu.rf_ram.memory[15][1] ;
 wire \u_cpu.rf_ram.memory[15][2] ;
 wire \u_cpu.rf_ram.memory[15][3] ;
 wire \u_cpu.rf_ram.memory[15][4] ;
 wire \u_cpu.rf_ram.memory[15][5] ;
 wire \u_cpu.rf_ram.memory[15][6] ;
 wire \u_cpu.rf_ram.memory[15][7] ;
 wire \u_cpu.rf_ram.memory[16][0] ;
 wire \u_cpu.rf_ram.memory[16][1] ;
 wire \u_cpu.rf_ram.memory[16][2] ;
 wire \u_cpu.rf_ram.memory[16][3] ;
 wire \u_cpu.rf_ram.memory[16][4] ;
 wire \u_cpu.rf_ram.memory[16][5] ;
 wire \u_cpu.rf_ram.memory[16][6] ;
 wire \u_cpu.rf_ram.memory[16][7] ;
 wire \u_cpu.rf_ram.memory[17][0] ;
 wire \u_cpu.rf_ram.memory[17][1] ;
 wire \u_cpu.rf_ram.memory[17][2] ;
 wire \u_cpu.rf_ram.memory[17][3] ;
 wire \u_cpu.rf_ram.memory[17][4] ;
 wire \u_cpu.rf_ram.memory[17][5] ;
 wire \u_cpu.rf_ram.memory[17][6] ;
 wire \u_cpu.rf_ram.memory[17][7] ;
 wire \u_cpu.rf_ram.memory[18][0] ;
 wire \u_cpu.rf_ram.memory[18][1] ;
 wire \u_cpu.rf_ram.memory[18][2] ;
 wire \u_cpu.rf_ram.memory[18][3] ;
 wire \u_cpu.rf_ram.memory[18][4] ;
 wire \u_cpu.rf_ram.memory[18][5] ;
 wire \u_cpu.rf_ram.memory[18][6] ;
 wire \u_cpu.rf_ram.memory[18][7] ;
 wire \u_cpu.rf_ram.memory[19][0] ;
 wire \u_cpu.rf_ram.memory[19][1] ;
 wire \u_cpu.rf_ram.memory[19][2] ;
 wire \u_cpu.rf_ram.memory[19][3] ;
 wire \u_cpu.rf_ram.memory[19][4] ;
 wire \u_cpu.rf_ram.memory[19][5] ;
 wire \u_cpu.rf_ram.memory[19][6] ;
 wire \u_cpu.rf_ram.memory[19][7] ;
 wire \u_cpu.rf_ram.memory[1][0] ;
 wire \u_cpu.rf_ram.memory[1][1] ;
 wire \u_cpu.rf_ram.memory[1][2] ;
 wire \u_cpu.rf_ram.memory[1][3] ;
 wire \u_cpu.rf_ram.memory[1][4] ;
 wire \u_cpu.rf_ram.memory[1][5] ;
 wire \u_cpu.rf_ram.memory[1][6] ;
 wire \u_cpu.rf_ram.memory[1][7] ;
 wire \u_cpu.rf_ram.memory[20][0] ;
 wire \u_cpu.rf_ram.memory[20][1] ;
 wire \u_cpu.rf_ram.memory[20][2] ;
 wire \u_cpu.rf_ram.memory[20][3] ;
 wire \u_cpu.rf_ram.memory[20][4] ;
 wire \u_cpu.rf_ram.memory[20][5] ;
 wire \u_cpu.rf_ram.memory[20][6] ;
 wire \u_cpu.rf_ram.memory[20][7] ;
 wire \u_cpu.rf_ram.memory[21][0] ;
 wire \u_cpu.rf_ram.memory[21][1] ;
 wire \u_cpu.rf_ram.memory[21][2] ;
 wire \u_cpu.rf_ram.memory[21][3] ;
 wire \u_cpu.rf_ram.memory[21][4] ;
 wire \u_cpu.rf_ram.memory[21][5] ;
 wire \u_cpu.rf_ram.memory[21][6] ;
 wire \u_cpu.rf_ram.memory[21][7] ;
 wire \u_cpu.rf_ram.memory[22][0] ;
 wire \u_cpu.rf_ram.memory[22][1] ;
 wire \u_cpu.rf_ram.memory[22][2] ;
 wire \u_cpu.rf_ram.memory[22][3] ;
 wire \u_cpu.rf_ram.memory[22][4] ;
 wire \u_cpu.rf_ram.memory[22][5] ;
 wire \u_cpu.rf_ram.memory[22][6] ;
 wire \u_cpu.rf_ram.memory[22][7] ;
 wire \u_cpu.rf_ram.memory[23][0] ;
 wire \u_cpu.rf_ram.memory[23][1] ;
 wire \u_cpu.rf_ram.memory[23][2] ;
 wire \u_cpu.rf_ram.memory[23][3] ;
 wire \u_cpu.rf_ram.memory[23][4] ;
 wire \u_cpu.rf_ram.memory[23][5] ;
 wire \u_cpu.rf_ram.memory[23][6] ;
 wire \u_cpu.rf_ram.memory[23][7] ;
 wire \u_cpu.rf_ram.memory[24][0] ;
 wire \u_cpu.rf_ram.memory[24][1] ;
 wire \u_cpu.rf_ram.memory[24][2] ;
 wire \u_cpu.rf_ram.memory[24][3] ;
 wire \u_cpu.rf_ram.memory[24][4] ;
 wire \u_cpu.rf_ram.memory[24][5] ;
 wire \u_cpu.rf_ram.memory[24][6] ;
 wire \u_cpu.rf_ram.memory[24][7] ;
 wire \u_cpu.rf_ram.memory[25][0] ;
 wire \u_cpu.rf_ram.memory[25][1] ;
 wire \u_cpu.rf_ram.memory[25][2] ;
 wire \u_cpu.rf_ram.memory[25][3] ;
 wire \u_cpu.rf_ram.memory[25][4] ;
 wire \u_cpu.rf_ram.memory[25][5] ;
 wire \u_cpu.rf_ram.memory[25][6] ;
 wire \u_cpu.rf_ram.memory[25][7] ;
 wire \u_cpu.rf_ram.memory[26][0] ;
 wire \u_cpu.rf_ram.memory[26][1] ;
 wire \u_cpu.rf_ram.memory[26][2] ;
 wire \u_cpu.rf_ram.memory[26][3] ;
 wire \u_cpu.rf_ram.memory[26][4] ;
 wire \u_cpu.rf_ram.memory[26][5] ;
 wire \u_cpu.rf_ram.memory[26][6] ;
 wire \u_cpu.rf_ram.memory[26][7] ;
 wire \u_cpu.rf_ram.memory[27][0] ;
 wire \u_cpu.rf_ram.memory[27][1] ;
 wire \u_cpu.rf_ram.memory[27][2] ;
 wire \u_cpu.rf_ram.memory[27][3] ;
 wire \u_cpu.rf_ram.memory[27][4] ;
 wire \u_cpu.rf_ram.memory[27][5] ;
 wire \u_cpu.rf_ram.memory[27][6] ;
 wire \u_cpu.rf_ram.memory[27][7] ;
 wire \u_cpu.rf_ram.memory[28][0] ;
 wire \u_cpu.rf_ram.memory[28][1] ;
 wire \u_cpu.rf_ram.memory[28][2] ;
 wire \u_cpu.rf_ram.memory[28][3] ;
 wire \u_cpu.rf_ram.memory[28][4] ;
 wire \u_cpu.rf_ram.memory[28][5] ;
 wire \u_cpu.rf_ram.memory[28][6] ;
 wire \u_cpu.rf_ram.memory[28][7] ;
 wire \u_cpu.rf_ram.memory[29][0] ;
 wire \u_cpu.rf_ram.memory[29][1] ;
 wire \u_cpu.rf_ram.memory[29][2] ;
 wire \u_cpu.rf_ram.memory[29][3] ;
 wire \u_cpu.rf_ram.memory[29][4] ;
 wire \u_cpu.rf_ram.memory[29][5] ;
 wire \u_cpu.rf_ram.memory[29][6] ;
 wire \u_cpu.rf_ram.memory[29][7] ;
 wire \u_cpu.rf_ram.memory[2][0] ;
 wire \u_cpu.rf_ram.memory[2][1] ;
 wire \u_cpu.rf_ram.memory[2][2] ;
 wire \u_cpu.rf_ram.memory[2][3] ;
 wire \u_cpu.rf_ram.memory[2][4] ;
 wire \u_cpu.rf_ram.memory[2][5] ;
 wire \u_cpu.rf_ram.memory[2][6] ;
 wire \u_cpu.rf_ram.memory[2][7] ;
 wire \u_cpu.rf_ram.memory[30][0] ;
 wire \u_cpu.rf_ram.memory[30][1] ;
 wire \u_cpu.rf_ram.memory[30][2] ;
 wire \u_cpu.rf_ram.memory[30][3] ;
 wire \u_cpu.rf_ram.memory[30][4] ;
 wire \u_cpu.rf_ram.memory[30][5] ;
 wire \u_cpu.rf_ram.memory[30][6] ;
 wire \u_cpu.rf_ram.memory[30][7] ;
 wire \u_cpu.rf_ram.memory[31][0] ;
 wire \u_cpu.rf_ram.memory[31][1] ;
 wire \u_cpu.rf_ram.memory[31][2] ;
 wire \u_cpu.rf_ram.memory[31][3] ;
 wire \u_cpu.rf_ram.memory[31][4] ;
 wire \u_cpu.rf_ram.memory[31][5] ;
 wire \u_cpu.rf_ram.memory[31][6] ;
 wire \u_cpu.rf_ram.memory[31][7] ;
 wire \u_cpu.rf_ram.memory[32][0] ;
 wire \u_cpu.rf_ram.memory[32][1] ;
 wire \u_cpu.rf_ram.memory[32][2] ;
 wire \u_cpu.rf_ram.memory[32][3] ;
 wire \u_cpu.rf_ram.memory[32][4] ;
 wire \u_cpu.rf_ram.memory[32][5] ;
 wire \u_cpu.rf_ram.memory[32][6] ;
 wire \u_cpu.rf_ram.memory[32][7] ;
 wire \u_cpu.rf_ram.memory[33][0] ;
 wire \u_cpu.rf_ram.memory[33][1] ;
 wire \u_cpu.rf_ram.memory[33][2] ;
 wire \u_cpu.rf_ram.memory[33][3] ;
 wire \u_cpu.rf_ram.memory[33][4] ;
 wire \u_cpu.rf_ram.memory[33][5] ;
 wire \u_cpu.rf_ram.memory[33][6] ;
 wire \u_cpu.rf_ram.memory[33][7] ;
 wire \u_cpu.rf_ram.memory[34][0] ;
 wire \u_cpu.rf_ram.memory[34][1] ;
 wire \u_cpu.rf_ram.memory[34][2] ;
 wire \u_cpu.rf_ram.memory[34][3] ;
 wire \u_cpu.rf_ram.memory[34][4] ;
 wire \u_cpu.rf_ram.memory[34][5] ;
 wire \u_cpu.rf_ram.memory[34][6] ;
 wire \u_cpu.rf_ram.memory[34][7] ;
 wire \u_cpu.rf_ram.memory[35][0] ;
 wire \u_cpu.rf_ram.memory[35][1] ;
 wire \u_cpu.rf_ram.memory[35][2] ;
 wire \u_cpu.rf_ram.memory[35][3] ;
 wire \u_cpu.rf_ram.memory[35][4] ;
 wire \u_cpu.rf_ram.memory[35][5] ;
 wire \u_cpu.rf_ram.memory[35][6] ;
 wire \u_cpu.rf_ram.memory[35][7] ;
 wire \u_cpu.rf_ram.memory[36][0] ;
 wire \u_cpu.rf_ram.memory[36][1] ;
 wire \u_cpu.rf_ram.memory[36][2] ;
 wire \u_cpu.rf_ram.memory[36][3] ;
 wire \u_cpu.rf_ram.memory[36][4] ;
 wire \u_cpu.rf_ram.memory[36][5] ;
 wire \u_cpu.rf_ram.memory[36][6] ;
 wire \u_cpu.rf_ram.memory[36][7] ;
 wire \u_cpu.rf_ram.memory[37][0] ;
 wire \u_cpu.rf_ram.memory[37][1] ;
 wire \u_cpu.rf_ram.memory[37][2] ;
 wire \u_cpu.rf_ram.memory[37][3] ;
 wire \u_cpu.rf_ram.memory[37][4] ;
 wire \u_cpu.rf_ram.memory[37][5] ;
 wire \u_cpu.rf_ram.memory[37][6] ;
 wire \u_cpu.rf_ram.memory[37][7] ;
 wire \u_cpu.rf_ram.memory[38][0] ;
 wire \u_cpu.rf_ram.memory[38][1] ;
 wire \u_cpu.rf_ram.memory[38][2] ;
 wire \u_cpu.rf_ram.memory[38][3] ;
 wire \u_cpu.rf_ram.memory[38][4] ;
 wire \u_cpu.rf_ram.memory[38][5] ;
 wire \u_cpu.rf_ram.memory[38][6] ;
 wire \u_cpu.rf_ram.memory[38][7] ;
 wire \u_cpu.rf_ram.memory[39][0] ;
 wire \u_cpu.rf_ram.memory[39][1] ;
 wire \u_cpu.rf_ram.memory[39][2] ;
 wire \u_cpu.rf_ram.memory[39][3] ;
 wire \u_cpu.rf_ram.memory[39][4] ;
 wire \u_cpu.rf_ram.memory[39][5] ;
 wire \u_cpu.rf_ram.memory[39][6] ;
 wire \u_cpu.rf_ram.memory[39][7] ;
 wire \u_cpu.rf_ram.memory[3][0] ;
 wire \u_cpu.rf_ram.memory[3][1] ;
 wire \u_cpu.rf_ram.memory[3][2] ;
 wire \u_cpu.rf_ram.memory[3][3] ;
 wire \u_cpu.rf_ram.memory[3][4] ;
 wire \u_cpu.rf_ram.memory[3][5] ;
 wire \u_cpu.rf_ram.memory[3][6] ;
 wire \u_cpu.rf_ram.memory[3][7] ;
 wire \u_cpu.rf_ram.memory[40][0] ;
 wire \u_cpu.rf_ram.memory[40][1] ;
 wire \u_cpu.rf_ram.memory[40][2] ;
 wire \u_cpu.rf_ram.memory[40][3] ;
 wire \u_cpu.rf_ram.memory[40][4] ;
 wire \u_cpu.rf_ram.memory[40][5] ;
 wire \u_cpu.rf_ram.memory[40][6] ;
 wire \u_cpu.rf_ram.memory[40][7] ;
 wire \u_cpu.rf_ram.memory[41][0] ;
 wire \u_cpu.rf_ram.memory[41][1] ;
 wire \u_cpu.rf_ram.memory[41][2] ;
 wire \u_cpu.rf_ram.memory[41][3] ;
 wire \u_cpu.rf_ram.memory[41][4] ;
 wire \u_cpu.rf_ram.memory[41][5] ;
 wire \u_cpu.rf_ram.memory[41][6] ;
 wire \u_cpu.rf_ram.memory[41][7] ;
 wire \u_cpu.rf_ram.memory[42][0] ;
 wire \u_cpu.rf_ram.memory[42][1] ;
 wire \u_cpu.rf_ram.memory[42][2] ;
 wire \u_cpu.rf_ram.memory[42][3] ;
 wire \u_cpu.rf_ram.memory[42][4] ;
 wire \u_cpu.rf_ram.memory[42][5] ;
 wire \u_cpu.rf_ram.memory[42][6] ;
 wire \u_cpu.rf_ram.memory[42][7] ;
 wire \u_cpu.rf_ram.memory[43][0] ;
 wire \u_cpu.rf_ram.memory[43][1] ;
 wire \u_cpu.rf_ram.memory[43][2] ;
 wire \u_cpu.rf_ram.memory[43][3] ;
 wire \u_cpu.rf_ram.memory[43][4] ;
 wire \u_cpu.rf_ram.memory[43][5] ;
 wire \u_cpu.rf_ram.memory[43][6] ;
 wire \u_cpu.rf_ram.memory[43][7] ;
 wire \u_cpu.rf_ram.memory[44][0] ;
 wire \u_cpu.rf_ram.memory[44][1] ;
 wire \u_cpu.rf_ram.memory[44][2] ;
 wire \u_cpu.rf_ram.memory[44][3] ;
 wire \u_cpu.rf_ram.memory[44][4] ;
 wire \u_cpu.rf_ram.memory[44][5] ;
 wire \u_cpu.rf_ram.memory[44][6] ;
 wire \u_cpu.rf_ram.memory[44][7] ;
 wire \u_cpu.rf_ram.memory[45][0] ;
 wire \u_cpu.rf_ram.memory[45][1] ;
 wire \u_cpu.rf_ram.memory[45][2] ;
 wire \u_cpu.rf_ram.memory[45][3] ;
 wire \u_cpu.rf_ram.memory[45][4] ;
 wire \u_cpu.rf_ram.memory[45][5] ;
 wire \u_cpu.rf_ram.memory[45][6] ;
 wire \u_cpu.rf_ram.memory[45][7] ;
 wire \u_cpu.rf_ram.memory[46][0] ;
 wire \u_cpu.rf_ram.memory[46][1] ;
 wire \u_cpu.rf_ram.memory[46][2] ;
 wire \u_cpu.rf_ram.memory[46][3] ;
 wire \u_cpu.rf_ram.memory[46][4] ;
 wire \u_cpu.rf_ram.memory[46][5] ;
 wire \u_cpu.rf_ram.memory[46][6] ;
 wire \u_cpu.rf_ram.memory[46][7] ;
 wire \u_cpu.rf_ram.memory[47][0] ;
 wire \u_cpu.rf_ram.memory[47][1] ;
 wire \u_cpu.rf_ram.memory[47][2] ;
 wire \u_cpu.rf_ram.memory[47][3] ;
 wire \u_cpu.rf_ram.memory[47][4] ;
 wire \u_cpu.rf_ram.memory[47][5] ;
 wire \u_cpu.rf_ram.memory[47][6] ;
 wire \u_cpu.rf_ram.memory[47][7] ;
 wire \u_cpu.rf_ram.memory[48][0] ;
 wire \u_cpu.rf_ram.memory[48][1] ;
 wire \u_cpu.rf_ram.memory[48][2] ;
 wire \u_cpu.rf_ram.memory[48][3] ;
 wire \u_cpu.rf_ram.memory[48][4] ;
 wire \u_cpu.rf_ram.memory[48][5] ;
 wire \u_cpu.rf_ram.memory[48][6] ;
 wire \u_cpu.rf_ram.memory[48][7] ;
 wire \u_cpu.rf_ram.memory[49][0] ;
 wire \u_cpu.rf_ram.memory[49][1] ;
 wire \u_cpu.rf_ram.memory[49][2] ;
 wire \u_cpu.rf_ram.memory[49][3] ;
 wire \u_cpu.rf_ram.memory[49][4] ;
 wire \u_cpu.rf_ram.memory[49][5] ;
 wire \u_cpu.rf_ram.memory[49][6] ;
 wire \u_cpu.rf_ram.memory[49][7] ;
 wire \u_cpu.rf_ram.memory[4][0] ;
 wire \u_cpu.rf_ram.memory[4][1] ;
 wire \u_cpu.rf_ram.memory[4][2] ;
 wire \u_cpu.rf_ram.memory[4][3] ;
 wire \u_cpu.rf_ram.memory[4][4] ;
 wire \u_cpu.rf_ram.memory[4][5] ;
 wire \u_cpu.rf_ram.memory[4][6] ;
 wire \u_cpu.rf_ram.memory[4][7] ;
 wire \u_cpu.rf_ram.memory[50][0] ;
 wire \u_cpu.rf_ram.memory[50][1] ;
 wire \u_cpu.rf_ram.memory[50][2] ;
 wire \u_cpu.rf_ram.memory[50][3] ;
 wire \u_cpu.rf_ram.memory[50][4] ;
 wire \u_cpu.rf_ram.memory[50][5] ;
 wire \u_cpu.rf_ram.memory[50][6] ;
 wire \u_cpu.rf_ram.memory[50][7] ;
 wire \u_cpu.rf_ram.memory[51][0] ;
 wire \u_cpu.rf_ram.memory[51][1] ;
 wire \u_cpu.rf_ram.memory[51][2] ;
 wire \u_cpu.rf_ram.memory[51][3] ;
 wire \u_cpu.rf_ram.memory[51][4] ;
 wire \u_cpu.rf_ram.memory[51][5] ;
 wire \u_cpu.rf_ram.memory[51][6] ;
 wire \u_cpu.rf_ram.memory[51][7] ;
 wire \u_cpu.rf_ram.memory[52][0] ;
 wire \u_cpu.rf_ram.memory[52][1] ;
 wire \u_cpu.rf_ram.memory[52][2] ;
 wire \u_cpu.rf_ram.memory[52][3] ;
 wire \u_cpu.rf_ram.memory[52][4] ;
 wire \u_cpu.rf_ram.memory[52][5] ;
 wire \u_cpu.rf_ram.memory[52][6] ;
 wire \u_cpu.rf_ram.memory[52][7] ;
 wire \u_cpu.rf_ram.memory[53][0] ;
 wire \u_cpu.rf_ram.memory[53][1] ;
 wire \u_cpu.rf_ram.memory[53][2] ;
 wire \u_cpu.rf_ram.memory[53][3] ;
 wire \u_cpu.rf_ram.memory[53][4] ;
 wire \u_cpu.rf_ram.memory[53][5] ;
 wire \u_cpu.rf_ram.memory[53][6] ;
 wire \u_cpu.rf_ram.memory[53][7] ;
 wire \u_cpu.rf_ram.memory[54][0] ;
 wire \u_cpu.rf_ram.memory[54][1] ;
 wire \u_cpu.rf_ram.memory[54][2] ;
 wire \u_cpu.rf_ram.memory[54][3] ;
 wire \u_cpu.rf_ram.memory[54][4] ;
 wire \u_cpu.rf_ram.memory[54][5] ;
 wire \u_cpu.rf_ram.memory[54][6] ;
 wire \u_cpu.rf_ram.memory[54][7] ;
 wire \u_cpu.rf_ram.memory[55][0] ;
 wire \u_cpu.rf_ram.memory[55][1] ;
 wire \u_cpu.rf_ram.memory[55][2] ;
 wire \u_cpu.rf_ram.memory[55][3] ;
 wire \u_cpu.rf_ram.memory[55][4] ;
 wire \u_cpu.rf_ram.memory[55][5] ;
 wire \u_cpu.rf_ram.memory[55][6] ;
 wire \u_cpu.rf_ram.memory[55][7] ;
 wire \u_cpu.rf_ram.memory[56][0] ;
 wire \u_cpu.rf_ram.memory[56][1] ;
 wire \u_cpu.rf_ram.memory[56][2] ;
 wire \u_cpu.rf_ram.memory[56][3] ;
 wire \u_cpu.rf_ram.memory[56][4] ;
 wire \u_cpu.rf_ram.memory[56][5] ;
 wire \u_cpu.rf_ram.memory[56][6] ;
 wire \u_cpu.rf_ram.memory[56][7] ;
 wire \u_cpu.rf_ram.memory[57][0] ;
 wire \u_cpu.rf_ram.memory[57][1] ;
 wire \u_cpu.rf_ram.memory[57][2] ;
 wire \u_cpu.rf_ram.memory[57][3] ;
 wire \u_cpu.rf_ram.memory[57][4] ;
 wire \u_cpu.rf_ram.memory[57][5] ;
 wire \u_cpu.rf_ram.memory[57][6] ;
 wire \u_cpu.rf_ram.memory[57][7] ;
 wire \u_cpu.rf_ram.memory[58][0] ;
 wire \u_cpu.rf_ram.memory[58][1] ;
 wire \u_cpu.rf_ram.memory[58][2] ;
 wire \u_cpu.rf_ram.memory[58][3] ;
 wire \u_cpu.rf_ram.memory[58][4] ;
 wire \u_cpu.rf_ram.memory[58][5] ;
 wire \u_cpu.rf_ram.memory[58][6] ;
 wire \u_cpu.rf_ram.memory[58][7] ;
 wire \u_cpu.rf_ram.memory[59][0] ;
 wire \u_cpu.rf_ram.memory[59][1] ;
 wire \u_cpu.rf_ram.memory[59][2] ;
 wire \u_cpu.rf_ram.memory[59][3] ;
 wire \u_cpu.rf_ram.memory[59][4] ;
 wire \u_cpu.rf_ram.memory[59][5] ;
 wire \u_cpu.rf_ram.memory[59][6] ;
 wire \u_cpu.rf_ram.memory[59][7] ;
 wire \u_cpu.rf_ram.memory[5][0] ;
 wire \u_cpu.rf_ram.memory[5][1] ;
 wire \u_cpu.rf_ram.memory[5][2] ;
 wire \u_cpu.rf_ram.memory[5][3] ;
 wire \u_cpu.rf_ram.memory[5][4] ;
 wire \u_cpu.rf_ram.memory[5][5] ;
 wire \u_cpu.rf_ram.memory[5][6] ;
 wire \u_cpu.rf_ram.memory[5][7] ;
 wire \u_cpu.rf_ram.memory[60][0] ;
 wire \u_cpu.rf_ram.memory[60][1] ;
 wire \u_cpu.rf_ram.memory[60][2] ;
 wire \u_cpu.rf_ram.memory[60][3] ;
 wire \u_cpu.rf_ram.memory[60][4] ;
 wire \u_cpu.rf_ram.memory[60][5] ;
 wire \u_cpu.rf_ram.memory[60][6] ;
 wire \u_cpu.rf_ram.memory[60][7] ;
 wire \u_cpu.rf_ram.memory[61][0] ;
 wire \u_cpu.rf_ram.memory[61][1] ;
 wire \u_cpu.rf_ram.memory[61][2] ;
 wire \u_cpu.rf_ram.memory[61][3] ;
 wire \u_cpu.rf_ram.memory[61][4] ;
 wire \u_cpu.rf_ram.memory[61][5] ;
 wire \u_cpu.rf_ram.memory[61][6] ;
 wire \u_cpu.rf_ram.memory[61][7] ;
 wire \u_cpu.rf_ram.memory[62][0] ;
 wire \u_cpu.rf_ram.memory[62][1] ;
 wire \u_cpu.rf_ram.memory[62][2] ;
 wire \u_cpu.rf_ram.memory[62][3] ;
 wire \u_cpu.rf_ram.memory[62][4] ;
 wire \u_cpu.rf_ram.memory[62][5] ;
 wire \u_cpu.rf_ram.memory[62][6] ;
 wire \u_cpu.rf_ram.memory[62][7] ;
 wire \u_cpu.rf_ram.memory[63][0] ;
 wire \u_cpu.rf_ram.memory[63][1] ;
 wire \u_cpu.rf_ram.memory[63][2] ;
 wire \u_cpu.rf_ram.memory[63][3] ;
 wire \u_cpu.rf_ram.memory[63][4] ;
 wire \u_cpu.rf_ram.memory[63][5] ;
 wire \u_cpu.rf_ram.memory[63][6] ;
 wire \u_cpu.rf_ram.memory[63][7] ;
 wire \u_cpu.rf_ram.memory[64][0] ;
 wire \u_cpu.rf_ram.memory[64][1] ;
 wire \u_cpu.rf_ram.memory[64][2] ;
 wire \u_cpu.rf_ram.memory[64][3] ;
 wire \u_cpu.rf_ram.memory[64][4] ;
 wire \u_cpu.rf_ram.memory[64][5] ;
 wire \u_cpu.rf_ram.memory[64][6] ;
 wire \u_cpu.rf_ram.memory[64][7] ;
 wire \u_cpu.rf_ram.memory[65][0] ;
 wire \u_cpu.rf_ram.memory[65][1] ;
 wire \u_cpu.rf_ram.memory[65][2] ;
 wire \u_cpu.rf_ram.memory[65][3] ;
 wire \u_cpu.rf_ram.memory[65][4] ;
 wire \u_cpu.rf_ram.memory[65][5] ;
 wire \u_cpu.rf_ram.memory[65][6] ;
 wire \u_cpu.rf_ram.memory[65][7] ;
 wire \u_cpu.rf_ram.memory[66][0] ;
 wire \u_cpu.rf_ram.memory[66][1] ;
 wire \u_cpu.rf_ram.memory[66][2] ;
 wire \u_cpu.rf_ram.memory[66][3] ;
 wire \u_cpu.rf_ram.memory[66][4] ;
 wire \u_cpu.rf_ram.memory[66][5] ;
 wire \u_cpu.rf_ram.memory[66][6] ;
 wire \u_cpu.rf_ram.memory[66][7] ;
 wire \u_cpu.rf_ram.memory[67][0] ;
 wire \u_cpu.rf_ram.memory[67][1] ;
 wire \u_cpu.rf_ram.memory[67][2] ;
 wire \u_cpu.rf_ram.memory[67][3] ;
 wire \u_cpu.rf_ram.memory[67][4] ;
 wire \u_cpu.rf_ram.memory[67][5] ;
 wire \u_cpu.rf_ram.memory[67][6] ;
 wire \u_cpu.rf_ram.memory[67][7] ;
 wire \u_cpu.rf_ram.memory[68][0] ;
 wire \u_cpu.rf_ram.memory[68][1] ;
 wire \u_cpu.rf_ram.memory[68][2] ;
 wire \u_cpu.rf_ram.memory[68][3] ;
 wire \u_cpu.rf_ram.memory[68][4] ;
 wire \u_cpu.rf_ram.memory[68][5] ;
 wire \u_cpu.rf_ram.memory[68][6] ;
 wire \u_cpu.rf_ram.memory[68][7] ;
 wire \u_cpu.rf_ram.memory[69][0] ;
 wire \u_cpu.rf_ram.memory[69][1] ;
 wire \u_cpu.rf_ram.memory[69][2] ;
 wire \u_cpu.rf_ram.memory[69][3] ;
 wire \u_cpu.rf_ram.memory[69][4] ;
 wire \u_cpu.rf_ram.memory[69][5] ;
 wire \u_cpu.rf_ram.memory[69][6] ;
 wire \u_cpu.rf_ram.memory[69][7] ;
 wire \u_cpu.rf_ram.memory[6][0] ;
 wire \u_cpu.rf_ram.memory[6][1] ;
 wire \u_cpu.rf_ram.memory[6][2] ;
 wire \u_cpu.rf_ram.memory[6][3] ;
 wire \u_cpu.rf_ram.memory[6][4] ;
 wire \u_cpu.rf_ram.memory[6][5] ;
 wire \u_cpu.rf_ram.memory[6][6] ;
 wire \u_cpu.rf_ram.memory[6][7] ;
 wire \u_cpu.rf_ram.memory[70][0] ;
 wire \u_cpu.rf_ram.memory[70][1] ;
 wire \u_cpu.rf_ram.memory[70][2] ;
 wire \u_cpu.rf_ram.memory[70][3] ;
 wire \u_cpu.rf_ram.memory[70][4] ;
 wire \u_cpu.rf_ram.memory[70][5] ;
 wire \u_cpu.rf_ram.memory[70][6] ;
 wire \u_cpu.rf_ram.memory[70][7] ;
 wire \u_cpu.rf_ram.memory[71][0] ;
 wire \u_cpu.rf_ram.memory[71][1] ;
 wire \u_cpu.rf_ram.memory[71][2] ;
 wire \u_cpu.rf_ram.memory[71][3] ;
 wire \u_cpu.rf_ram.memory[71][4] ;
 wire \u_cpu.rf_ram.memory[71][5] ;
 wire \u_cpu.rf_ram.memory[71][6] ;
 wire \u_cpu.rf_ram.memory[71][7] ;
 wire \u_cpu.rf_ram.memory[72][0] ;
 wire \u_cpu.rf_ram.memory[72][1] ;
 wire \u_cpu.rf_ram.memory[72][2] ;
 wire \u_cpu.rf_ram.memory[72][3] ;
 wire \u_cpu.rf_ram.memory[72][4] ;
 wire \u_cpu.rf_ram.memory[72][5] ;
 wire \u_cpu.rf_ram.memory[72][6] ;
 wire \u_cpu.rf_ram.memory[72][7] ;
 wire \u_cpu.rf_ram.memory[73][0] ;
 wire \u_cpu.rf_ram.memory[73][1] ;
 wire \u_cpu.rf_ram.memory[73][2] ;
 wire \u_cpu.rf_ram.memory[73][3] ;
 wire \u_cpu.rf_ram.memory[73][4] ;
 wire \u_cpu.rf_ram.memory[73][5] ;
 wire \u_cpu.rf_ram.memory[73][6] ;
 wire \u_cpu.rf_ram.memory[73][7] ;
 wire \u_cpu.rf_ram.memory[74][0] ;
 wire \u_cpu.rf_ram.memory[74][1] ;
 wire \u_cpu.rf_ram.memory[74][2] ;
 wire \u_cpu.rf_ram.memory[74][3] ;
 wire \u_cpu.rf_ram.memory[74][4] ;
 wire \u_cpu.rf_ram.memory[74][5] ;
 wire \u_cpu.rf_ram.memory[74][6] ;
 wire \u_cpu.rf_ram.memory[74][7] ;
 wire \u_cpu.rf_ram.memory[75][0] ;
 wire \u_cpu.rf_ram.memory[75][1] ;
 wire \u_cpu.rf_ram.memory[75][2] ;
 wire \u_cpu.rf_ram.memory[75][3] ;
 wire \u_cpu.rf_ram.memory[75][4] ;
 wire \u_cpu.rf_ram.memory[75][5] ;
 wire \u_cpu.rf_ram.memory[75][6] ;
 wire \u_cpu.rf_ram.memory[75][7] ;
 wire \u_cpu.rf_ram.memory[76][0] ;
 wire \u_cpu.rf_ram.memory[76][1] ;
 wire \u_cpu.rf_ram.memory[76][2] ;
 wire \u_cpu.rf_ram.memory[76][3] ;
 wire \u_cpu.rf_ram.memory[76][4] ;
 wire \u_cpu.rf_ram.memory[76][5] ;
 wire \u_cpu.rf_ram.memory[76][6] ;
 wire \u_cpu.rf_ram.memory[76][7] ;
 wire \u_cpu.rf_ram.memory[77][0] ;
 wire \u_cpu.rf_ram.memory[77][1] ;
 wire \u_cpu.rf_ram.memory[77][2] ;
 wire \u_cpu.rf_ram.memory[77][3] ;
 wire \u_cpu.rf_ram.memory[77][4] ;
 wire \u_cpu.rf_ram.memory[77][5] ;
 wire \u_cpu.rf_ram.memory[77][6] ;
 wire \u_cpu.rf_ram.memory[77][7] ;
 wire \u_cpu.rf_ram.memory[78][0] ;
 wire \u_cpu.rf_ram.memory[78][1] ;
 wire \u_cpu.rf_ram.memory[78][2] ;
 wire \u_cpu.rf_ram.memory[78][3] ;
 wire \u_cpu.rf_ram.memory[78][4] ;
 wire \u_cpu.rf_ram.memory[78][5] ;
 wire \u_cpu.rf_ram.memory[78][6] ;
 wire \u_cpu.rf_ram.memory[78][7] ;
 wire \u_cpu.rf_ram.memory[79][0] ;
 wire \u_cpu.rf_ram.memory[79][1] ;
 wire \u_cpu.rf_ram.memory[79][2] ;
 wire \u_cpu.rf_ram.memory[79][3] ;
 wire \u_cpu.rf_ram.memory[79][4] ;
 wire \u_cpu.rf_ram.memory[79][5] ;
 wire \u_cpu.rf_ram.memory[79][6] ;
 wire \u_cpu.rf_ram.memory[79][7] ;
 wire \u_cpu.rf_ram.memory[7][0] ;
 wire \u_cpu.rf_ram.memory[7][1] ;
 wire \u_cpu.rf_ram.memory[7][2] ;
 wire \u_cpu.rf_ram.memory[7][3] ;
 wire \u_cpu.rf_ram.memory[7][4] ;
 wire \u_cpu.rf_ram.memory[7][5] ;
 wire \u_cpu.rf_ram.memory[7][6] ;
 wire \u_cpu.rf_ram.memory[7][7] ;
 wire \u_cpu.rf_ram.memory[80][0] ;
 wire \u_cpu.rf_ram.memory[80][1] ;
 wire \u_cpu.rf_ram.memory[80][2] ;
 wire \u_cpu.rf_ram.memory[80][3] ;
 wire \u_cpu.rf_ram.memory[80][4] ;
 wire \u_cpu.rf_ram.memory[80][5] ;
 wire \u_cpu.rf_ram.memory[80][6] ;
 wire \u_cpu.rf_ram.memory[80][7] ;
 wire \u_cpu.rf_ram.memory[81][0] ;
 wire \u_cpu.rf_ram.memory[81][1] ;
 wire \u_cpu.rf_ram.memory[81][2] ;
 wire \u_cpu.rf_ram.memory[81][3] ;
 wire \u_cpu.rf_ram.memory[81][4] ;
 wire \u_cpu.rf_ram.memory[81][5] ;
 wire \u_cpu.rf_ram.memory[81][6] ;
 wire \u_cpu.rf_ram.memory[81][7] ;
 wire \u_cpu.rf_ram.memory[82][0] ;
 wire \u_cpu.rf_ram.memory[82][1] ;
 wire \u_cpu.rf_ram.memory[82][2] ;
 wire \u_cpu.rf_ram.memory[82][3] ;
 wire \u_cpu.rf_ram.memory[82][4] ;
 wire \u_cpu.rf_ram.memory[82][5] ;
 wire \u_cpu.rf_ram.memory[82][6] ;
 wire \u_cpu.rf_ram.memory[82][7] ;
 wire \u_cpu.rf_ram.memory[83][0] ;
 wire \u_cpu.rf_ram.memory[83][1] ;
 wire \u_cpu.rf_ram.memory[83][2] ;
 wire \u_cpu.rf_ram.memory[83][3] ;
 wire \u_cpu.rf_ram.memory[83][4] ;
 wire \u_cpu.rf_ram.memory[83][5] ;
 wire \u_cpu.rf_ram.memory[83][6] ;
 wire \u_cpu.rf_ram.memory[83][7] ;
 wire \u_cpu.rf_ram.memory[84][0] ;
 wire \u_cpu.rf_ram.memory[84][1] ;
 wire \u_cpu.rf_ram.memory[84][2] ;
 wire \u_cpu.rf_ram.memory[84][3] ;
 wire \u_cpu.rf_ram.memory[84][4] ;
 wire \u_cpu.rf_ram.memory[84][5] ;
 wire \u_cpu.rf_ram.memory[84][6] ;
 wire \u_cpu.rf_ram.memory[84][7] ;
 wire \u_cpu.rf_ram.memory[85][0] ;
 wire \u_cpu.rf_ram.memory[85][1] ;
 wire \u_cpu.rf_ram.memory[85][2] ;
 wire \u_cpu.rf_ram.memory[85][3] ;
 wire \u_cpu.rf_ram.memory[85][4] ;
 wire \u_cpu.rf_ram.memory[85][5] ;
 wire \u_cpu.rf_ram.memory[85][6] ;
 wire \u_cpu.rf_ram.memory[85][7] ;
 wire \u_cpu.rf_ram.memory[86][0] ;
 wire \u_cpu.rf_ram.memory[86][1] ;
 wire \u_cpu.rf_ram.memory[86][2] ;
 wire \u_cpu.rf_ram.memory[86][3] ;
 wire \u_cpu.rf_ram.memory[86][4] ;
 wire \u_cpu.rf_ram.memory[86][5] ;
 wire \u_cpu.rf_ram.memory[86][6] ;
 wire \u_cpu.rf_ram.memory[86][7] ;
 wire \u_cpu.rf_ram.memory[87][0] ;
 wire \u_cpu.rf_ram.memory[87][1] ;
 wire \u_cpu.rf_ram.memory[87][2] ;
 wire \u_cpu.rf_ram.memory[87][3] ;
 wire \u_cpu.rf_ram.memory[87][4] ;
 wire \u_cpu.rf_ram.memory[87][5] ;
 wire \u_cpu.rf_ram.memory[87][6] ;
 wire \u_cpu.rf_ram.memory[87][7] ;
 wire \u_cpu.rf_ram.memory[88][0] ;
 wire \u_cpu.rf_ram.memory[88][1] ;
 wire \u_cpu.rf_ram.memory[88][2] ;
 wire \u_cpu.rf_ram.memory[88][3] ;
 wire \u_cpu.rf_ram.memory[88][4] ;
 wire \u_cpu.rf_ram.memory[88][5] ;
 wire \u_cpu.rf_ram.memory[88][6] ;
 wire \u_cpu.rf_ram.memory[88][7] ;
 wire \u_cpu.rf_ram.memory[89][0] ;
 wire \u_cpu.rf_ram.memory[89][1] ;
 wire \u_cpu.rf_ram.memory[89][2] ;
 wire \u_cpu.rf_ram.memory[89][3] ;
 wire \u_cpu.rf_ram.memory[89][4] ;
 wire \u_cpu.rf_ram.memory[89][5] ;
 wire \u_cpu.rf_ram.memory[89][6] ;
 wire \u_cpu.rf_ram.memory[89][7] ;
 wire \u_cpu.rf_ram.memory[8][0] ;
 wire \u_cpu.rf_ram.memory[8][1] ;
 wire \u_cpu.rf_ram.memory[8][2] ;
 wire \u_cpu.rf_ram.memory[8][3] ;
 wire \u_cpu.rf_ram.memory[8][4] ;
 wire \u_cpu.rf_ram.memory[8][5] ;
 wire \u_cpu.rf_ram.memory[8][6] ;
 wire \u_cpu.rf_ram.memory[8][7] ;
 wire \u_cpu.rf_ram.memory[90][0] ;
 wire \u_cpu.rf_ram.memory[90][1] ;
 wire \u_cpu.rf_ram.memory[90][2] ;
 wire \u_cpu.rf_ram.memory[90][3] ;
 wire \u_cpu.rf_ram.memory[90][4] ;
 wire \u_cpu.rf_ram.memory[90][5] ;
 wire \u_cpu.rf_ram.memory[90][6] ;
 wire \u_cpu.rf_ram.memory[90][7] ;
 wire \u_cpu.rf_ram.memory[91][0] ;
 wire \u_cpu.rf_ram.memory[91][1] ;
 wire \u_cpu.rf_ram.memory[91][2] ;
 wire \u_cpu.rf_ram.memory[91][3] ;
 wire \u_cpu.rf_ram.memory[91][4] ;
 wire \u_cpu.rf_ram.memory[91][5] ;
 wire \u_cpu.rf_ram.memory[91][6] ;
 wire \u_cpu.rf_ram.memory[91][7] ;
 wire \u_cpu.rf_ram.memory[92][0] ;
 wire \u_cpu.rf_ram.memory[92][1] ;
 wire \u_cpu.rf_ram.memory[92][2] ;
 wire \u_cpu.rf_ram.memory[92][3] ;
 wire \u_cpu.rf_ram.memory[92][4] ;
 wire \u_cpu.rf_ram.memory[92][5] ;
 wire \u_cpu.rf_ram.memory[92][6] ;
 wire \u_cpu.rf_ram.memory[92][7] ;
 wire \u_cpu.rf_ram.memory[93][0] ;
 wire \u_cpu.rf_ram.memory[93][1] ;
 wire \u_cpu.rf_ram.memory[93][2] ;
 wire \u_cpu.rf_ram.memory[93][3] ;
 wire \u_cpu.rf_ram.memory[93][4] ;
 wire \u_cpu.rf_ram.memory[93][5] ;
 wire \u_cpu.rf_ram.memory[93][6] ;
 wire \u_cpu.rf_ram.memory[93][7] ;
 wire \u_cpu.rf_ram.memory[94][0] ;
 wire \u_cpu.rf_ram.memory[94][1] ;
 wire \u_cpu.rf_ram.memory[94][2] ;
 wire \u_cpu.rf_ram.memory[94][3] ;
 wire \u_cpu.rf_ram.memory[94][4] ;
 wire \u_cpu.rf_ram.memory[94][5] ;
 wire \u_cpu.rf_ram.memory[94][6] ;
 wire \u_cpu.rf_ram.memory[94][7] ;
 wire \u_cpu.rf_ram.memory[95][0] ;
 wire \u_cpu.rf_ram.memory[95][1] ;
 wire \u_cpu.rf_ram.memory[95][2] ;
 wire \u_cpu.rf_ram.memory[95][3] ;
 wire \u_cpu.rf_ram.memory[95][4] ;
 wire \u_cpu.rf_ram.memory[95][5] ;
 wire \u_cpu.rf_ram.memory[95][6] ;
 wire \u_cpu.rf_ram.memory[95][7] ;
 wire \u_cpu.rf_ram.memory[96][0] ;
 wire \u_cpu.rf_ram.memory[96][1] ;
 wire \u_cpu.rf_ram.memory[96][2] ;
 wire \u_cpu.rf_ram.memory[96][3] ;
 wire \u_cpu.rf_ram.memory[96][4] ;
 wire \u_cpu.rf_ram.memory[96][5] ;
 wire \u_cpu.rf_ram.memory[96][6] ;
 wire \u_cpu.rf_ram.memory[96][7] ;
 wire \u_cpu.rf_ram.memory[97][0] ;
 wire \u_cpu.rf_ram.memory[97][1] ;
 wire \u_cpu.rf_ram.memory[97][2] ;
 wire \u_cpu.rf_ram.memory[97][3] ;
 wire \u_cpu.rf_ram.memory[97][4] ;
 wire \u_cpu.rf_ram.memory[97][5] ;
 wire \u_cpu.rf_ram.memory[97][6] ;
 wire \u_cpu.rf_ram.memory[97][7] ;
 wire \u_cpu.rf_ram.memory[98][0] ;
 wire \u_cpu.rf_ram.memory[98][1] ;
 wire \u_cpu.rf_ram.memory[98][2] ;
 wire \u_cpu.rf_ram.memory[98][3] ;
 wire \u_cpu.rf_ram.memory[98][4] ;
 wire \u_cpu.rf_ram.memory[98][5] ;
 wire \u_cpu.rf_ram.memory[98][6] ;
 wire \u_cpu.rf_ram.memory[98][7] ;
 wire \u_cpu.rf_ram.memory[99][0] ;
 wire \u_cpu.rf_ram.memory[99][1] ;
 wire \u_cpu.rf_ram.memory[99][2] ;
 wire \u_cpu.rf_ram.memory[99][3] ;
 wire \u_cpu.rf_ram.memory[99][4] ;
 wire \u_cpu.rf_ram.memory[99][5] ;
 wire \u_cpu.rf_ram.memory[99][6] ;
 wire \u_cpu.rf_ram.memory[99][7] ;
 wire \u_cpu.rf_ram.memory[9][0] ;
 wire \u_cpu.rf_ram.memory[9][1] ;
 wire \u_cpu.rf_ram.memory[9][2] ;
 wire \u_cpu.rf_ram.memory[9][3] ;
 wire \u_cpu.rf_ram.memory[9][4] ;
 wire \u_cpu.rf_ram.memory[9][5] ;
 wire \u_cpu.rf_ram.memory[9][6] ;
 wire \u_cpu.rf_ram.memory[9][7] ;
 wire \u_cpu.rf_ram.rdata[0] ;
 wire \u_cpu.rf_ram.rdata[1] ;
 wire \u_cpu.rf_ram.rdata[2] ;
 wire \u_cpu.rf_ram.rdata[3] ;
 wire \u_cpu.rf_ram.rdata[4] ;
 wire \u_cpu.rf_ram.rdata[5] ;
 wire \u_cpu.rf_ram.rdata[6] ;
 wire \u_cpu.rf_ram.rdata[7] ;
 wire \u_cpu.rf_ram.regzero ;
 wire \u_cpu.rf_ram_if.genblk1.wtrig0_r ;
 wire \u_cpu.rf_ram_if.rcnt[0] ;
 wire \u_cpu.rf_ram_if.rcnt[1] ;
 wire \u_cpu.rf_ram_if.rcnt[2] ;
 wire \u_cpu.rf_ram_if.rdata0[1] ;
 wire \u_cpu.rf_ram_if.rdata0[2] ;
 wire \u_cpu.rf_ram_if.rdata0[3] ;
 wire \u_cpu.rf_ram_if.rdata0[4] ;
 wire \u_cpu.rf_ram_if.rdata0[5] ;
 wire \u_cpu.rf_ram_if.rdata0[6] ;
 wire \u_cpu.rf_ram_if.rdata0[7] ;
 wire \u_cpu.rf_ram_if.rdata1[0] ;
 wire \u_cpu.rf_ram_if.rdata1[1] ;
 wire \u_cpu.rf_ram_if.rdata1[2] ;
 wire \u_cpu.rf_ram_if.rdata1[3] ;
 wire \u_cpu.rf_ram_if.rdata1[4] ;
 wire \u_cpu.rf_ram_if.rdata1[5] ;
 wire \u_cpu.rf_ram_if.rdata1[6] ;
 wire \u_cpu.rf_ram_if.rgnt ;
 wire \u_cpu.rf_ram_if.rreq_r ;
 wire \u_cpu.rf_ram_if.rtrig0 ;
 wire \u_cpu.rf_ram_if.rtrig1 ;
 wire \u_cpu.rf_ram_if.wdata0_r[0] ;
 wire \u_cpu.rf_ram_if.wdata0_r[1] ;
 wire \u_cpu.rf_ram_if.wdata0_r[2] ;
 wire \u_cpu.rf_ram_if.wdata0_r[3] ;
 wire \u_cpu.rf_ram_if.wdata0_r[4] ;
 wire \u_cpu.rf_ram_if.wdata0_r[5] ;
 wire \u_cpu.rf_ram_if.wdata0_r[6] ;
 wire \u_cpu.rf_ram_if.wdata1_r[0] ;
 wire \u_cpu.rf_ram_if.wdata1_r[1] ;
 wire \u_cpu.rf_ram_if.wdata1_r[2] ;
 wire \u_cpu.rf_ram_if.wdata1_r[3] ;
 wire \u_cpu.rf_ram_if.wdata1_r[4] ;
 wire \u_cpu.rf_ram_if.wdata1_r[5] ;
 wire \u_cpu.rf_ram_if.wdata1_r[6] ;
 wire \u_cpu.rf_ram_if.wdata1_r[7] ;
 wire \u_cpu.rf_ram_if.wen0_r ;
 wire \u_cpu.rf_ram_if.wen1_r ;
 wire \u_cpu.rf_ram_if.wtrig0 ;
 wire \u_scanchain_local.clk ;
 wire \u_scanchain_local.clk_out ;
 wire \u_scanchain_local.data_out ;
 wire \u_scanchain_local.data_out_i ;
 wire \u_scanchain_local.module_data_in[34] ;
 wire \u_scanchain_local.module_data_in[35] ;
 wire \u_scanchain_local.module_data_in[36] ;
 wire \u_scanchain_local.module_data_in[37] ;
 wire \u_scanchain_local.module_data_in[38] ;
 wire \u_scanchain_local.module_data_in[39] ;
 wire \u_scanchain_local.module_data_in[40] ;
 wire \u_scanchain_local.module_data_in[41] ;
 wire \u_scanchain_local.module_data_in[42] ;
 wire \u_scanchain_local.module_data_in[43] ;
 wire \u_scanchain_local.module_data_in[44] ;
 wire \u_scanchain_local.module_data_in[45] ;
 wire \u_scanchain_local.module_data_in[46] ;
 wire \u_scanchain_local.module_data_in[47] ;
 wire \u_scanchain_local.module_data_in[48] ;
 wire \u_scanchain_local.module_data_in[49] ;
 wire \u_scanchain_local.module_data_in[50] ;
 wire \u_scanchain_local.module_data_in[51] ;
 wire \u_scanchain_local.module_data_in[52] ;
 wire \u_scanchain_local.module_data_in[53] ;
 wire \u_scanchain_local.module_data_in[54] ;
 wire \u_scanchain_local.module_data_in[55] ;
 wire \u_scanchain_local.module_data_in[56] ;
 wire \u_scanchain_local.module_data_in[57] ;
 wire \u_scanchain_local.module_data_in[58] ;
 wire \u_scanchain_local.module_data_in[59] ;
 wire \u_scanchain_local.module_data_in[60] ;
 wire \u_scanchain_local.module_data_in[61] ;
 wire \u_scanchain_local.module_data_in[62] ;
 wire \u_scanchain_local.module_data_in[63] ;
 wire \u_scanchain_local.module_data_in[64] ;
 wire \u_scanchain_local.module_data_in[65] ;
 wire \u_scanchain_local.module_data_in[66] ;
 wire \u_scanchain_local.module_data_in[67] ;
 wire \u_scanchain_local.module_data_in[68] ;
 wire \u_scanchain_local.module_data_in[69] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;

 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05713_ (.I(\u_cpu.rf_ram_if.rcnt[0] ),
    .ZN(_01366_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _05714_ (.A1(\u_cpu.rf_ram_if.rcnt[2] ),
    .A2(\u_cpu.rf_ram_if.rcnt[1] ),
    .A3(_01366_),
    .Z(_01367_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05715_ (.I(_01367_),
    .ZN(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05716_ (.I(_01368_),
    .Z(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05717_ (.I(\u_cpu.cpu.bufreg.lsb[0] ),
    .Z(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05718_ (.I(\u_cpu.cpu.bufreg.lsb[1] ),
    .Z(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05719_ (.A1(_01369_),
    .A2(_01370_),
    .ZN(\u_arbiter.i_wb_cpu_dbus_sel[0] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05720_ (.I(\u_cpu.cpu.decode.co_mem_word ),
    .Z(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05721_ (.I(\u_cpu.cpu.bne_or_bge ),
    .Z(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _05722_ (.A1(\u_cpu.cpu.csr_d_sel ),
    .A2(_01371_),
    .A3(_01372_),
    .ZN(_01373_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05723_ (.I(\u_cpu.cpu.decode.opcode[2] ),
    .Z(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05724_ (.I(_01374_),
    .ZN(_01375_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05725_ (.I(\u_cpu.cpu.branch_op ),
    .ZN(_01376_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05726_ (.A1(_01375_),
    .A2(_01376_),
    .ZN(_01377_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _05727_ (.A1(\u_cpu.cpu.decode.op21 ),
    .A2(_01373_),
    .A3(_01377_),
    .ZN(_01378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _05728_ (.A1(\u_cpu.cpu.decode.opcode[2] ),
    .A2(\u_cpu.cpu.branch_op ),
    .ZN(_01379_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05729_ (.A1(_01373_),
    .A2(_01379_),
    .ZN(_01380_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05730_ (.I(\u_cpu.cpu.decode.op26 ),
    .ZN(_01381_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05731_ (.I(\u_cpu.cpu.decode.co_ebreak ),
    .ZN(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05732_ (.A1(\u_cpu.cpu.decode.op21 ),
    .A2(_01381_),
    .B(_01382_),
    .ZN(_01383_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _05733_ (.A1(\u_cpu.cpu.csr_d_sel ),
    .A2(\u_cpu.cpu.decode.co_mem_word ),
    .A3(\u_cpu.cpu.decode.op21 ),
    .A4(_01372_),
    .Z(_01384_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05734_ (.I(\u_cpu.cpu.genblk3.csr.o_new_irq ),
    .ZN(_01385_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05735_ (.I(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ),
    .ZN(_01386_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _05736_ (.A1(_01379_),
    .A2(_01384_),
    .B(_01385_),
    .C(_01386_),
    .ZN(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _05737_ (.A1(_01380_),
    .A2(_01383_),
    .B(_01387_),
    .ZN(_01388_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _05738_ (.A1(_01368_),
    .A2(_01378_),
    .A3(_01388_),
    .Z(_01389_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05739_ (.A1(\u_cpu.cpu.immdec.imm24_20[0] ),
    .A2(_01389_),
    .Z(_01390_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05740_ (.I(\u_cpu.cpu.csr_imm ),
    .ZN(_01391_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05741_ (.A1(_01391_),
    .A2(_01368_),
    .ZN(_01392_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05742_ (.A1(_01379_),
    .A2(_01384_),
    .ZN(_01393_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _05743_ (.A1(\u_cpu.cpu.genblk3.csr.o_new_irq ),
    .A2(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ),
    .A3(_01393_),
    .ZN(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05744_ (.A1(\u_cpu.cpu.decode.op21 ),
    .A2(_01381_),
    .ZN(_01395_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _05745_ (.A1(_01394_),
    .A2(_01395_),
    .B(_01388_),
    .C(_01367_),
    .ZN(_01396_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _05746_ (.A1(_01390_),
    .A2(_01392_),
    .A3(_01396_),
    .Z(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05747_ (.I(_01397_),
    .Z(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05748_ (.I(_01398_),
    .Z(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05749_ (.I(_01399_),
    .Z(_01400_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05750_ (.I(_01367_),
    .Z(_01401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05751_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[8] ),
    .A2(_01401_),
    .ZN(_01402_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05752_ (.A1(\u_cpu.cpu.immdec.imm24_20[4] ),
    .A2(_01389_),
    .ZN(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05753_ (.A1(_01402_),
    .A2(_01403_),
    .ZN(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _05754_ (.A1(_01378_),
    .A2(_01388_),
    .B(_01401_),
    .ZN(_01405_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05755_ (.A1(_01404_),
    .A2(_01405_),
    .ZN(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05756_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[5] ),
    .A2(\u_cpu.rf_ram_if.rtrig0 ),
    .ZN(_01407_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05757_ (.I(\u_cpu.cpu.csr_d_sel ),
    .Z(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05758_ (.I(_01408_),
    .ZN(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05759_ (.A1(\u_cpu.cpu.decode.co_mem_word ),
    .A2(\u_cpu.cpu.bne_or_bge ),
    .ZN(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05760_ (.I(_01410_),
    .Z(_01411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05761_ (.A1(_01409_),
    .A2(_01411_),
    .ZN(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05762_ (.A1(_01412_),
    .A2(_01377_),
    .ZN(_01413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05763_ (.A1(\u_cpu.cpu.decode.op26 ),
    .A2(\u_cpu.cpu.decode.co_ebreak ),
    .ZN(_01414_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _05764_ (.A1(_01413_),
    .A2(_01414_),
    .B(\u_cpu.rf_ram_if.rtrig0 ),
    .C(_01378_),
    .ZN(_01415_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05765_ (.A1(\u_cpu.cpu.immdec.imm24_20[1] ),
    .A2(_01388_),
    .B(_01415_),
    .ZN(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05766_ (.A1(_01407_),
    .A2(_01416_),
    .Z(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05767_ (.I(_01417_),
    .Z(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05768_ (.I(_01418_),
    .Z(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05769_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[7] ),
    .A2(_01367_),
    .ZN(_01420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05770_ (.A1(\u_cpu.cpu.immdec.imm24_20[3] ),
    .A2(_01389_),
    .ZN(_01421_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05771_ (.A1(_01420_),
    .A2(_01421_),
    .Z(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05772_ (.I(_01422_),
    .Z(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05773_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[6] ),
    .A2(_01367_),
    .ZN(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05774_ (.A1(\u_cpu.cpu.immdec.imm24_20[2] ),
    .A2(_01389_),
    .ZN(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05775_ (.A1(_01424_),
    .A2(_01425_),
    .Z(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05776_ (.I(_01426_),
    .Z(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05777_ (.I(_01427_),
    .Z(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _05778_ (.A1(_01406_),
    .A2(_01419_),
    .A3(_01423_),
    .A4(_01428_),
    .ZN(_01429_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05779_ (.A1(_01400_),
    .A2(_01429_),
    .ZN(_00025_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05780_ (.I(_01401_),
    .Z(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05781_ (.I(_01430_),
    .ZN(\u_cpu.rf_ram_if.wtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05782_ (.I(\u_arbiter.i_wb_cpu_ibus_adr[0] ),
    .Z(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05783_ (.I(net2),
    .ZN(_01432_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05784_ (.A1(_01432_),
    .A2(\u_cpu.cpu.state.ibus_cyc ),
    .Z(_01433_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05785_ (.I(_01433_),
    .Z(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05786_ (.A1(_01431_),
    .A2(_01434_),
    .Z(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05787_ (.I(_01435_),
    .Z(\u_arbiter.o_wb_cpu_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05788_ (.A1(\u_arbiter.i_wb_cpu_ibus_adr[1] ),
    .A2(_01433_),
    .Z(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05789_ (.I(_01436_),
    .Z(\u_arbiter.o_wb_cpu_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05790_ (.I(\u_cpu.cpu.genblk1.align.ctrl_misal ),
    .Z(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05791_ (.I(_01437_),
    .Z(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05792_ (.I(_01438_),
    .Z(_01439_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05793_ (.I(_01439_),
    .Z(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05794_ (.I(_01440_),
    .Z(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05795_ (.I(_01441_),
    .Z(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05796_ (.I(_01442_),
    .Z(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05797_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[2] ),
    .Z(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05798_ (.A1(_01443_),
    .A2(_01444_),
    .ZN(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05799_ (.I(_01441_),
    .Z(_01446_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05800_ (.I(_01446_),
    .Z(_01447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05801_ (.A1(_01447_),
    .A2(_01444_),
    .ZN(_01448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05802_ (.A1(_01434_),
    .A2(_01448_),
    .ZN(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05803_ (.A1(_01432_),
    .A2(\u_cpu.cpu.state.ibus_cyc ),
    .ZN(_01450_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05804_ (.I(_01450_),
    .Z(_01451_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05805_ (.I(_01451_),
    .Z(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05806_ (.I(_01452_),
    .Z(_01453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05807_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[2] ),
    .A2(_01453_),
    .ZN(_01454_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05808_ (.A1(_01445_),
    .A2(_01449_),
    .B(_01454_),
    .ZN(\u_arbiter.o_wb_cpu_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05809_ (.I(_01451_),
    .Z(_01455_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05810_ (.I(_01455_),
    .Z(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05811_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[3] ),
    .A2(_01448_),
    .Z(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05812_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[3] ),
    .A2(_01453_),
    .ZN(_01458_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05813_ (.A1(_01456_),
    .A2(_01457_),
    .B(_01458_),
    .ZN(\u_arbiter.o_wb_cpu_adr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05814_ (.A1(_01447_),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[3] ),
    .A3(_01444_),
    .ZN(_01459_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05815_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[4] ),
    .A2(_01459_),
    .Z(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05816_ (.I(_01452_),
    .Z(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05817_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[4] ),
    .A2(_01461_),
    .ZN(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05818_ (.A1(_01456_),
    .A2(_01460_),
    .B(_01462_),
    .ZN(\u_arbiter.o_wb_cpu_adr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05819_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[5] ),
    .Z(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _05820_ (.A1(\u_cpu.cpu.genblk1.align.ctrl_misal ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[4] ),
    .A3(\u_cpu.cpu.ctrl.o_ibus_adr[3] ),
    .A4(\u_cpu.cpu.ctrl.o_ibus_adr[2] ),
    .Z(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05821_ (.A1(_01463_),
    .A2(_01464_),
    .ZN(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05822_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[5] ),
    .A2(_01461_),
    .ZN(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05823_ (.A1(_01456_),
    .A2(_01465_),
    .B(_01466_),
    .ZN(\u_arbiter.o_wb_cpu_adr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05824_ (.A1(_01463_),
    .A2(_01464_),
    .B(\u_cpu.cpu.ctrl.o_ibus_adr[6] ),
    .ZN(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05825_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[6] ),
    .A2(_01463_),
    .A3(_01464_),
    .ZN(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05826_ (.A1(_01434_),
    .A2(_01468_),
    .ZN(_01469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05827_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[6] ),
    .A2(_01461_),
    .ZN(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05828_ (.A1(_01467_),
    .A2(_01469_),
    .B(_01470_),
    .ZN(\u_arbiter.o_wb_cpu_adr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05829_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[7] ),
    .A2(_01468_),
    .Z(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05830_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[7] ),
    .A2(_01461_),
    .ZN(_01472_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05831_ (.A1(_01456_),
    .A2(_01471_),
    .B(_01472_),
    .ZN(\u_arbiter.o_wb_cpu_adr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05832_ (.I(_01455_),
    .Z(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05833_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[8] ),
    .ZN(_01474_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _05834_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[7] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[6] ),
    .A3(\u_cpu.cpu.ctrl.o_ibus_adr[5] ),
    .A4(_01464_),
    .ZN(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05835_ (.A1(_01474_),
    .A2(_01475_),
    .ZN(_01476_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05836_ (.A1(_01474_),
    .A2(_01475_),
    .Z(_01477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05837_ (.A1(_01476_),
    .A2(_01477_),
    .ZN(_01478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05838_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[8] ),
    .A2(_01461_),
    .ZN(_01479_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05839_ (.A1(_01473_),
    .A2(_01478_),
    .B(_01479_),
    .ZN(\u_arbiter.o_wb_cpu_adr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05840_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[9] ),
    .A2(_01477_),
    .Z(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05841_ (.I(_01452_),
    .Z(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05842_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[9] ),
    .A2(_01481_),
    .ZN(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05843_ (.A1(_01473_),
    .A2(_01480_),
    .B(_01482_),
    .ZN(\u_arbiter.o_wb_cpu_adr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05844_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[10] ),
    .A2(_01453_),
    .ZN(_01483_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05845_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[10] ),
    .Z(_01484_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05846_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[9] ),
    .ZN(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05847_ (.A1(_01485_),
    .A2(_01477_),
    .ZN(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05848_ (.A1(_01484_),
    .A2(_01486_),
    .B(_01455_),
    .ZN(_01487_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05849_ (.A1(_01484_),
    .A2(_01486_),
    .B(_01487_),
    .ZN(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05850_ (.A1(_01483_),
    .A2(_01488_),
    .ZN(\u_arbiter.o_wb_cpu_adr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05851_ (.I(_01452_),
    .Z(_01489_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05852_ (.A1(_01484_),
    .A2(_01486_),
    .B(\u_cpu.cpu.ctrl.o_ibus_adr[11] ),
    .ZN(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05853_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[11] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[10] ),
    .ZN(_01491_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _05854_ (.A1(_01485_),
    .A2(_01474_),
    .A3(_01475_),
    .A4(_01491_),
    .ZN(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05855_ (.I(_01451_),
    .Z(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05856_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[11] ),
    .A2(_01493_),
    .ZN(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05857_ (.A1(_01489_),
    .A2(_01490_),
    .A3(_01492_),
    .B(_01494_),
    .ZN(\u_arbiter.o_wb_cpu_adr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05858_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[12] ),
    .Z(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05859_ (.A1(_01495_),
    .A2(_01492_),
    .ZN(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05860_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[12] ),
    .A2(_01481_),
    .ZN(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05861_ (.A1(_01473_),
    .A2(_01496_),
    .B(_01497_),
    .ZN(\u_arbiter.o_wb_cpu_adr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05862_ (.A1(_01495_),
    .A2(_01492_),
    .B(\u_cpu.cpu.ctrl.o_ibus_adr[13] ),
    .ZN(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _05863_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[13] ),
    .A2(_01495_),
    .A3(_01492_),
    .Z(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05864_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[13] ),
    .A2(_01493_),
    .ZN(_01500_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05865_ (.A1(_01489_),
    .A2(_01498_),
    .A3(_01499_),
    .B(_01500_),
    .ZN(\u_arbiter.o_wb_cpu_adr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05866_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[14] ),
    .A2(_01453_),
    .ZN(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05867_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[14] ),
    .Z(_01502_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05868_ (.A1(_01502_),
    .A2(_01499_),
    .B(_01455_),
    .ZN(_01503_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05869_ (.A1(_01502_),
    .A2(_01499_),
    .B(_01503_),
    .ZN(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05870_ (.A1(_01501_),
    .A2(_01504_),
    .ZN(\u_arbiter.o_wb_cpu_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05871_ (.I(_01452_),
    .Z(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05872_ (.A1(_01502_),
    .A2(_01499_),
    .B(\u_cpu.cpu.ctrl.o_ibus_adr[15] ),
    .ZN(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05873_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[15] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[14] ),
    .Z(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _05874_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[13] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[12] ),
    .A3(_01492_),
    .A4(_01507_),
    .Z(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05875_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[15] ),
    .A2(_01493_),
    .ZN(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05876_ (.A1(_01505_),
    .A2(_01506_),
    .A3(_01508_),
    .B(_01509_),
    .ZN(\u_arbiter.o_wb_cpu_adr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05877_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[16] ),
    .A2(_01508_),
    .ZN(_01510_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05878_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[16] ),
    .A2(_01508_),
    .Z(_01511_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05879_ (.I(_01451_),
    .Z(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05880_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[16] ),
    .A2(_01512_),
    .ZN(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05881_ (.A1(_01505_),
    .A2(_01510_),
    .A3(_01511_),
    .B(_01513_),
    .ZN(\u_arbiter.o_wb_cpu_adr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05882_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[17] ),
    .A2(_01511_),
    .ZN(_01514_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05883_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[17] ),
    .A2(_01481_),
    .ZN(_01515_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05884_ (.A1(_01473_),
    .A2(_01514_),
    .B(_01515_),
    .ZN(\u_arbiter.o_wb_cpu_adr[17] ));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _05885_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[18] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[17] ),
    .A3(\u_cpu.cpu.ctrl.o_ibus_adr[16] ),
    .A4(_01508_),
    .Z(_01516_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05886_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[17] ),
    .A2(_01511_),
    .B(\u_cpu.cpu.ctrl.o_ibus_adr[18] ),
    .ZN(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05887_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[18] ),
    .A2(_01512_),
    .ZN(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05888_ (.A1(_01505_),
    .A2(_01516_),
    .A3(_01517_),
    .B(_01518_),
    .ZN(\u_arbiter.o_wb_cpu_adr[18] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05889_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[19] ),
    .A2(_01516_),
    .Z(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05890_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[19] ),
    .A2(_01516_),
    .ZN(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05891_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[19] ),
    .A2(_01512_),
    .ZN(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05892_ (.A1(_01505_),
    .A2(_01519_),
    .A3(_01520_),
    .B(_01521_),
    .ZN(\u_arbiter.o_wb_cpu_adr[19] ));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05893_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[20] ),
    .A2(_01519_),
    .ZN(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05894_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[20] ),
    .A2(_01481_),
    .ZN(_01523_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05895_ (.A1(_01473_),
    .A2(_01522_),
    .B(_01523_),
    .ZN(\u_arbiter.o_wb_cpu_adr[20] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05896_ (.I(_01455_),
    .Z(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05897_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[20] ),
    .A2(_01519_),
    .ZN(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05898_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[21] ),
    .A2(_01525_),
    .Z(_01526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05899_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[21] ),
    .A2(_01481_),
    .ZN(_01527_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05900_ (.A1(_01524_),
    .A2(_01526_),
    .B(_01527_),
    .ZN(\u_arbiter.o_wb_cpu_adr[21] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05901_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[22] ),
    .ZN(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _05902_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[21] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[20] ),
    .A3(\u_cpu.cpu.ctrl.o_ibus_adr[19] ),
    .A4(_01516_),
    .ZN(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05903_ (.A1(_01528_),
    .A2(_01529_),
    .Z(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05904_ (.A1(_01528_),
    .A2(_01529_),
    .ZN(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05905_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[22] ),
    .A2(_01512_),
    .ZN(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05906_ (.A1(_01505_),
    .A2(_01530_),
    .A3(_01531_),
    .B(_01532_),
    .ZN(\u_arbiter.o_wb_cpu_adr[22] ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05907_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[23] ),
    .A2(_01531_),
    .ZN(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05908_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[23] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[22] ),
    .ZN(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05909_ (.A1(_01529_),
    .A2(_01534_),
    .ZN(_01535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05910_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[23] ),
    .A2(_01512_),
    .ZN(_01536_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05911_ (.A1(_01453_),
    .A2(_01533_),
    .A3(_01535_),
    .B(_01536_),
    .ZN(\u_arbiter.o_wb_cpu_adr[23] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05912_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[24] ),
    .Z(_01537_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05913_ (.A1(_01537_),
    .A2(_01535_),
    .ZN(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05914_ (.I(_01451_),
    .Z(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05915_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[24] ),
    .A2(_01539_),
    .ZN(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05916_ (.A1(_01524_),
    .A2(_01538_),
    .B(_01540_),
    .ZN(\u_arbiter.o_wb_cpu_adr[24] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05917_ (.A1(_01537_),
    .A2(_01535_),
    .ZN(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05918_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[25] ),
    .A2(_01541_),
    .Z(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05919_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[25] ),
    .A2(_01539_),
    .ZN(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05920_ (.A1(_01524_),
    .A2(_01542_),
    .B(_01543_),
    .ZN(\u_arbiter.o_wb_cpu_adr[25] ));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05921_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[25] ),
    .A2(_01537_),
    .A3(_01535_),
    .ZN(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05922_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[26] ),
    .A2(_01544_),
    .Z(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05923_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[26] ),
    .A2(_01539_),
    .ZN(_01546_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05924_ (.A1(_01524_),
    .A2(_01545_),
    .B(_01546_),
    .ZN(\u_arbiter.o_wb_cpu_adr[26] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05925_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[27] ),
    .Z(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _05926_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[26] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[25] ),
    .A3(\u_cpu.cpu.ctrl.o_ibus_adr[24] ),
    .A4(_01535_),
    .Z(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05927_ (.A1(_01547_),
    .A2(_01548_),
    .ZN(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05928_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[27] ),
    .A2(_01539_),
    .ZN(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05929_ (.A1(_01524_),
    .A2(_01549_),
    .B(_01550_),
    .ZN(\u_arbiter.o_wb_cpu_adr[27] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05930_ (.A1(_01547_),
    .A2(_01548_),
    .ZN(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05931_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[28] ),
    .A2(_01551_),
    .Z(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05932_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[28] ),
    .A2(_01539_),
    .ZN(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05933_ (.A1(_01489_),
    .A2(_01552_),
    .B(_01553_),
    .ZN(\u_arbiter.o_wb_cpu_adr[28] ));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05934_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[28] ),
    .A2(_01547_),
    .A3(_01548_),
    .ZN(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05935_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[29] ),
    .A2(_01554_),
    .Z(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05936_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[29] ),
    .A2(_01493_),
    .ZN(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05937_ (.A1(_01489_),
    .A2(_01555_),
    .B(_01556_),
    .ZN(\u_arbiter.o_wb_cpu_adr[29] ));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _05938_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[29] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[28] ),
    .A3(\u_cpu.cpu.ctrl.o_ibus_adr[27] ),
    .A4(_01548_),
    .ZN(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05939_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[30] ),
    .A2(_01557_),
    .Z(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05940_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[30] ),
    .A2(_01493_),
    .ZN(_01559_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05941_ (.A1(_01489_),
    .A2(_01558_),
    .B(_01559_),
    .ZN(\u_arbiter.o_wb_cpu_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05942_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[30] ),
    .ZN(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05943_ (.A1(_01560_),
    .A2(_01557_),
    .ZN(_01561_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05944_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[31] ),
    .A2(_01561_),
    .Z(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05945_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[31] ),
    .I1(_01562_),
    .S(_01434_),
    .Z(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05946_ (.I(_01563_),
    .Z(\u_arbiter.o_wb_cpu_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05947_ (.I(_01406_),
    .Z(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05948_ (.A1(_01420_),
    .A2(_01421_),
    .ZN(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05949_ (.I(_01565_),
    .Z(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _05950_ (.A1(_01390_),
    .A2(_01392_),
    .A3(_01396_),
    .ZN(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05951_ (.I(_01567_),
    .Z(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05952_ (.I(_01568_),
    .Z(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05953_ (.I(_01569_),
    .Z(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05954_ (.I(\u_cpu.raddr[0] ),
    .Z(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05955_ (.I(_01571_),
    .Z(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05956_ (.I(_01572_),
    .Z(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05957_ (.I(_01573_),
    .Z(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05958_ (.I(\u_cpu.raddr[1] ),
    .Z(_01575_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05959_ (.I(_01575_),
    .Z(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05960_ (.I(_01576_),
    .Z(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05961_ (.I0(\u_cpu.rf_ram.memory[8][0] ),
    .I1(\u_cpu.rf_ram.memory[9][0] ),
    .I2(\u_cpu.rf_ram.memory[10][0] ),
    .I3(\u_cpu.rf_ram.memory[11][0] ),
    .S0(_01574_),
    .S1(_01577_),
    .Z(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05962_ (.A1(_01570_),
    .A2(_01578_),
    .ZN(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05963_ (.I(_01398_),
    .Z(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05964_ (.I(\u_cpu.raddr[0] ),
    .Z(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05965_ (.I(_01581_),
    .Z(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05966_ (.I(_01582_),
    .Z(_01583_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05967_ (.I(_01575_),
    .Z(_01584_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05968_ (.I(_01584_),
    .Z(_01585_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05969_ (.I0(\u_cpu.rf_ram.memory[12][0] ),
    .I1(\u_cpu.rf_ram.memory[13][0] ),
    .I2(\u_cpu.rf_ram.memory[14][0] ),
    .I3(\u_cpu.rf_ram.memory[15][0] ),
    .S0(_01583_),
    .S1(_01585_),
    .Z(_01586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05970_ (.I(_01417_),
    .Z(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05971_ (.I(_01587_),
    .Z(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05972_ (.A1(_01580_),
    .A2(_01586_),
    .B(_01588_),
    .ZN(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05973_ (.I(_01398_),
    .Z(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05974_ (.I(_01573_),
    .Z(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05975_ (.I(_01576_),
    .Z(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05976_ (.I0(\u_cpu.rf_ram.memory[4][0] ),
    .I1(\u_cpu.rf_ram.memory[5][0] ),
    .I2(\u_cpu.rf_ram.memory[6][0] ),
    .I3(\u_cpu.rf_ram.memory[7][0] ),
    .S0(_01591_),
    .S1(_01592_),
    .Z(_01593_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05977_ (.A1(_01590_),
    .A2(_01593_),
    .ZN(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05978_ (.I(_01567_),
    .Z(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05979_ (.I(_01595_),
    .Z(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05980_ (.I(_01596_),
    .Z(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05981_ (.I(_01582_),
    .Z(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05982_ (.I(_01584_),
    .Z(_01599_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05983_ (.I0(\u_cpu.rf_ram.memory[0][0] ),
    .I1(\u_cpu.rf_ram.memory[1][0] ),
    .I2(\u_cpu.rf_ram.memory[2][0] ),
    .I3(\u_cpu.rf_ram.memory[3][0] ),
    .S0(_01598_),
    .S1(_01599_),
    .Z(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05984_ (.A1(_01407_),
    .A2(_01416_),
    .ZN(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05985_ (.I(_01601_),
    .Z(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05986_ (.I(_01602_),
    .Z(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05987_ (.A1(_01597_),
    .A2(_01600_),
    .B(_01603_),
    .ZN(_01604_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05988_ (.A1(_01424_),
    .A2(_01425_),
    .ZN(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05989_ (.I(_01605_),
    .Z(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05990_ (.I(_01606_),
    .Z(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _05991_ (.A1(_01579_),
    .A2(_01589_),
    .B1(_01594_),
    .B2(_01604_),
    .C(_01607_),
    .ZN(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05992_ (.I(_01397_),
    .Z(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05993_ (.I(_01609_),
    .Z(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05994_ (.I(_01610_),
    .Z(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05995_ (.I(_01581_),
    .Z(_01612_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05996_ (.I(_01612_),
    .Z(_01613_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05997_ (.I(_01613_),
    .Z(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05998_ (.I(_01575_),
    .Z(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05999_ (.I(_01615_),
    .Z(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06000_ (.I0(\u_cpu.rf_ram.memory[20][0] ),
    .I1(\u_cpu.rf_ram.memory[21][0] ),
    .I2(\u_cpu.rf_ram.memory[22][0] ),
    .I3(\u_cpu.rf_ram.memory[23][0] ),
    .S0(_01614_),
    .S1(_01616_),
    .Z(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06001_ (.A1(_01611_),
    .A2(_01617_),
    .ZN(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06002_ (.I(_01596_),
    .Z(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06003_ (.I(_01571_),
    .Z(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06004_ (.I(_01620_),
    .Z(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06005_ (.I(_01621_),
    .Z(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06006_ (.I(\u_cpu.raddr[1] ),
    .Z(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06007_ (.I(_01623_),
    .Z(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06008_ (.I(_01624_),
    .Z(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06009_ (.I0(\u_cpu.rf_ram.memory[16][0] ),
    .I1(\u_cpu.rf_ram.memory[17][0] ),
    .I2(\u_cpu.rf_ram.memory[18][0] ),
    .I3(\u_cpu.rf_ram.memory[19][0] ),
    .S0(_01622_),
    .S1(_01625_),
    .Z(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06010_ (.I(_01601_),
    .Z(_01627_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06011_ (.I(_01627_),
    .Z(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06012_ (.A1(_01619_),
    .A2(_01626_),
    .B(_01628_),
    .ZN(_01629_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06013_ (.I(_01398_),
    .Z(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06014_ (.I(_01573_),
    .Z(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06015_ (.I(_01623_),
    .Z(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06016_ (.I(_01632_),
    .Z(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06017_ (.I(_01633_),
    .Z(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06018_ (.I0(\u_cpu.rf_ram.memory[28][0] ),
    .I1(\u_cpu.rf_ram.memory[29][0] ),
    .I2(\u_cpu.rf_ram.memory[30][0] ),
    .I3(\u_cpu.rf_ram.memory[31][0] ),
    .S0(_01631_),
    .S1(_01634_),
    .Z(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06019_ (.A1(_01630_),
    .A2(_01635_),
    .ZN(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06020_ (.I(_01596_),
    .Z(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06021_ (.I(_01571_),
    .Z(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06022_ (.I(_01638_),
    .Z(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06023_ (.I(_01639_),
    .Z(_01640_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06024_ (.I(_01575_),
    .Z(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06025_ (.I(_01641_),
    .Z(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06026_ (.I0(\u_cpu.rf_ram.memory[24][0] ),
    .I1(\u_cpu.rf_ram.memory[25][0] ),
    .I2(\u_cpu.rf_ram.memory[26][0] ),
    .I3(\u_cpu.rf_ram.memory[27][0] ),
    .S0(_01640_),
    .S1(_01642_),
    .Z(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06027_ (.I(_01418_),
    .Z(_01644_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06028_ (.A1(_01637_),
    .A2(_01643_),
    .B(_01644_),
    .ZN(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06029_ (.A1(_01618_),
    .A2(_01629_),
    .B1(_01636_),
    .B2(_01645_),
    .C(_01428_),
    .ZN(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06030_ (.I(_01422_),
    .Z(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06031_ (.I(_01397_),
    .Z(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06032_ (.I(_01648_),
    .Z(_01649_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06033_ (.I(_01581_),
    .Z(_01650_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06034_ (.I(_01650_),
    .Z(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06035_ (.I(_01623_),
    .Z(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06036_ (.I(_01652_),
    .Z(_01653_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06037_ (.I0(\u_cpu.rf_ram.memory[52][0] ),
    .I1(\u_cpu.rf_ram.memory[53][0] ),
    .I2(\u_cpu.rf_ram.memory[54][0] ),
    .I3(\u_cpu.rf_ram.memory[55][0] ),
    .S0(_01651_),
    .S1(_01653_),
    .Z(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06038_ (.A1(_01649_),
    .A2(_01654_),
    .ZN(_01655_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06039_ (.I(_01595_),
    .Z(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06040_ (.I(_01620_),
    .Z(_01657_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06041_ (.I(\u_cpu.raddr[1] ),
    .Z(_01658_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06042_ (.I(_01658_),
    .Z(_01659_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06043_ (.I(_01659_),
    .Z(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06044_ (.I0(\u_cpu.rf_ram.memory[48][0] ),
    .I1(\u_cpu.rf_ram.memory[49][0] ),
    .I2(\u_cpu.rf_ram.memory[50][0] ),
    .I3(\u_cpu.rf_ram.memory[51][0] ),
    .S0(_01657_),
    .S1(_01660_),
    .Z(_01661_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06045_ (.I(_01601_),
    .Z(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06046_ (.I(_01662_),
    .Z(_01663_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06047_ (.A1(_01656_),
    .A2(_01661_),
    .B(_01663_),
    .ZN(_01664_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06048_ (.I(_01397_),
    .Z(_01665_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06049_ (.I(_01665_),
    .Z(_01666_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06050_ (.I(_01623_),
    .Z(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06051_ (.I(_01667_),
    .Z(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06052_ (.I0(\u_cpu.rf_ram.memory[60][0] ),
    .I1(\u_cpu.rf_ram.memory[61][0] ),
    .I2(\u_cpu.rf_ram.memory[62][0] ),
    .I3(\u_cpu.rf_ram.memory[63][0] ),
    .S0(_01639_),
    .S1(_01668_),
    .Z(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06053_ (.A1(_01666_),
    .A2(_01669_),
    .ZN(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06054_ (.I(_01567_),
    .Z(_01671_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06055_ (.I(_01671_),
    .Z(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06056_ (.I(_01571_),
    .Z(_01673_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06057_ (.I(_01673_),
    .Z(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06058_ (.I(_01658_),
    .Z(_01675_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06059_ (.I(_01675_),
    .Z(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06060_ (.I0(\u_cpu.rf_ram.memory[56][0] ),
    .I1(\u_cpu.rf_ram.memory[57][0] ),
    .I2(\u_cpu.rf_ram.memory[58][0] ),
    .I3(\u_cpu.rf_ram.memory[59][0] ),
    .S0(_01674_),
    .S1(_01676_),
    .Z(_01677_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06061_ (.I(_01417_),
    .Z(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06062_ (.I(_01678_),
    .Z(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06063_ (.A1(_01672_),
    .A2(_01677_),
    .B(_01679_),
    .ZN(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06064_ (.I(_01426_),
    .Z(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06065_ (.A1(_01655_),
    .A2(_01664_),
    .B1(_01670_),
    .B2(_01680_),
    .C(_01681_),
    .ZN(_01682_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06066_ (.I(_01568_),
    .Z(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06067_ (.I(_01683_),
    .Z(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06068_ (.I(_01581_),
    .Z(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06069_ (.I(_01685_),
    .Z(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06070_ (.I(_01623_),
    .Z(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06071_ (.I(_01687_),
    .Z(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06072_ (.I0(\u_cpu.rf_ram.memory[40][0] ),
    .I1(\u_cpu.rf_ram.memory[41][0] ),
    .I2(\u_cpu.rf_ram.memory[42][0] ),
    .I3(\u_cpu.rf_ram.memory[43][0] ),
    .S0(_01686_),
    .S1(_01688_),
    .Z(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06073_ (.A1(_01684_),
    .A2(_01689_),
    .ZN(_01690_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06074_ (.I(_01609_),
    .Z(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06075_ (.I(_01620_),
    .Z(_01692_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06076_ (.I(_01659_),
    .Z(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06077_ (.I0(\u_cpu.rf_ram.memory[44][0] ),
    .I1(\u_cpu.rf_ram.memory[45][0] ),
    .I2(\u_cpu.rf_ram.memory[46][0] ),
    .I3(\u_cpu.rf_ram.memory[47][0] ),
    .S0(_01692_),
    .S1(_01693_),
    .Z(_01694_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06078_ (.I(_01678_),
    .Z(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06079_ (.A1(_01691_),
    .A2(_01694_),
    .B(_01695_),
    .ZN(_01696_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06080_ (.I(_01648_),
    .Z(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06081_ (.I(_01650_),
    .Z(_01698_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06082_ (.I(_01667_),
    .Z(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06083_ (.I0(\u_cpu.rf_ram.memory[36][0] ),
    .I1(\u_cpu.rf_ram.memory[37][0] ),
    .I2(\u_cpu.rf_ram.memory[38][0] ),
    .I3(\u_cpu.rf_ram.memory[39][0] ),
    .S0(_01698_),
    .S1(_01699_),
    .Z(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06084_ (.A1(_01697_),
    .A2(_01700_),
    .ZN(_01701_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06085_ (.I(_01567_),
    .Z(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06086_ (.I(_01702_),
    .Z(_01703_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06087_ (.I(_01571_),
    .Z(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06088_ (.I(_01704_),
    .Z(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06089_ (.I(_01658_),
    .Z(_01706_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06090_ (.I(_01706_),
    .Z(_01707_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06091_ (.I0(\u_cpu.rf_ram.memory[32][0] ),
    .I1(\u_cpu.rf_ram.memory[33][0] ),
    .I2(\u_cpu.rf_ram.memory[34][0] ),
    .I3(\u_cpu.rf_ram.memory[35][0] ),
    .S0(_01705_),
    .S1(_01707_),
    .Z(_01708_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06092_ (.I(_01662_),
    .Z(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06093_ (.A1(_01703_),
    .A2(_01708_),
    .B(_01709_),
    .ZN(_01710_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06094_ (.I(_01605_),
    .Z(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06095_ (.A1(_01690_),
    .A2(_01696_),
    .B1(_01701_),
    .B2(_01710_),
    .C(_01711_),
    .ZN(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06096_ (.A1(_01647_),
    .A2(_01682_),
    .A3(_01712_),
    .Z(_01713_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06097_ (.A1(_01566_),
    .A2(_01608_),
    .A3(_01646_),
    .B(_01713_),
    .ZN(_01714_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06098_ (.I(_01665_),
    .Z(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06099_ (.I(_01638_),
    .Z(_01716_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06100_ (.I(_01667_),
    .Z(_01717_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06101_ (.I0(\u_cpu.rf_ram.memory[108][0] ),
    .I1(\u_cpu.rf_ram.memory[109][0] ),
    .I2(\u_cpu.rf_ram.memory[110][0] ),
    .I3(\u_cpu.rf_ram.memory[111][0] ),
    .S0(_01716_),
    .S1(_01717_),
    .Z(_01718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06102_ (.A1(_01715_),
    .A2(_01718_),
    .ZN(_01719_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06103_ (.I(_01595_),
    .Z(_01720_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06104_ (.I(_01620_),
    .Z(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06105_ (.I0(\u_cpu.rf_ram.memory[104][0] ),
    .I1(\u_cpu.rf_ram.memory[105][0] ),
    .I2(\u_cpu.rf_ram.memory[106][0] ),
    .I3(\u_cpu.rf_ram.memory[107][0] ),
    .S0(_01721_),
    .S1(_01624_),
    .Z(_01722_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06106_ (.I(_01417_),
    .Z(_01723_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06107_ (.A1(_01720_),
    .A2(_01722_),
    .B(_01723_),
    .ZN(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06108_ (.I(_01665_),
    .Z(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06109_ (.I0(\u_cpu.rf_ram.memory[100][0] ),
    .I1(\u_cpu.rf_ram.memory[101][0] ),
    .I2(\u_cpu.rf_ram.memory[102][0] ),
    .I3(\u_cpu.rf_ram.memory[103][0] ),
    .S0(_01621_),
    .S1(_01633_),
    .Z(_01726_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06110_ (.A1(_01725_),
    .A2(_01726_),
    .ZN(_01727_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06111_ (.I(_01595_),
    .Z(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06112_ (.I(_01673_),
    .Z(_01729_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06113_ (.I0(\u_cpu.rf_ram.memory[96][0] ),
    .I1(\u_cpu.rf_ram.memory[97][0] ),
    .I2(\u_cpu.rf_ram.memory[98][0] ),
    .I3(\u_cpu.rf_ram.memory[99][0] ),
    .S0(_01729_),
    .S1(_01641_),
    .Z(_01730_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06114_ (.I(_01662_),
    .Z(_01731_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06115_ (.A1(_01728_),
    .A2(_01730_),
    .B(_01731_),
    .ZN(_01732_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06116_ (.I(_01605_),
    .Z(_01733_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06117_ (.A1(_01719_),
    .A2(_01724_),
    .B1(_01727_),
    .B2(_01732_),
    .C(_01733_),
    .ZN(_01734_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06118_ (.I(_01648_),
    .Z(_01735_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06119_ (.I(_01685_),
    .Z(_01736_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06120_ (.I(_01687_),
    .Z(_01737_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06121_ (.I0(\u_cpu.rf_ram.memory[124][0] ),
    .I1(\u_cpu.rf_ram.memory[125][0] ),
    .I2(\u_cpu.rf_ram.memory[126][0] ),
    .I3(\u_cpu.rf_ram.memory[127][0] ),
    .S0(_01736_),
    .S1(_01737_),
    .Z(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06122_ (.A1(_01735_),
    .A2(_01738_),
    .ZN(_01739_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06123_ (.I(_01671_),
    .Z(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06124_ (.I(_01673_),
    .Z(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06125_ (.I(_01675_),
    .Z(_01742_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06126_ (.I0(\u_cpu.rf_ram.memory[120][0] ),
    .I1(\u_cpu.rf_ram.memory[121][0] ),
    .I2(\u_cpu.rf_ram.memory[122][0] ),
    .I3(\u_cpu.rf_ram.memory[123][0] ),
    .S0(_01741_),
    .S1(_01742_),
    .Z(_01743_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06127_ (.I(_01678_),
    .Z(_01744_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06128_ (.A1(_01740_),
    .A2(_01743_),
    .B(_01744_),
    .ZN(_01745_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06129_ (.I(_01702_),
    .Z(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06130_ (.I(_01650_),
    .Z(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06131_ (.I(_01652_),
    .Z(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06132_ (.I0(\u_cpu.rf_ram.memory[112][0] ),
    .I1(\u_cpu.rf_ram.memory[113][0] ),
    .I2(\u_cpu.rf_ram.memory[114][0] ),
    .I3(\u_cpu.rf_ram.memory[115][0] ),
    .S0(_01747_),
    .S1(_01748_),
    .Z(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06133_ (.A1(_01746_),
    .A2(_01749_),
    .ZN(_01750_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06134_ (.I(_01609_),
    .Z(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06135_ (.I(_01704_),
    .Z(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06136_ (.I(_01706_),
    .Z(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06137_ (.I0(\u_cpu.rf_ram.memory[116][0] ),
    .I1(\u_cpu.rf_ram.memory[117][0] ),
    .I2(\u_cpu.rf_ram.memory[118][0] ),
    .I3(\u_cpu.rf_ram.memory[119][0] ),
    .S0(_01752_),
    .S1(_01753_),
    .Z(_01754_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06138_ (.I(_01662_),
    .Z(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06139_ (.A1(_01751_),
    .A2(_01754_),
    .B(_01755_),
    .ZN(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06140_ (.I(_01426_),
    .Z(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06141_ (.A1(_01739_),
    .A2(_01745_),
    .B1(_01750_),
    .B2(_01756_),
    .C(_01757_),
    .ZN(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06142_ (.A1(_01423_),
    .A2(_01734_),
    .A3(_01758_),
    .ZN(_01759_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06143_ (.I(_01565_),
    .Z(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06144_ (.I(_01648_),
    .Z(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06145_ (.I(_01612_),
    .Z(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06146_ (.I(_01687_),
    .Z(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06147_ (.I0(\u_cpu.rf_ram.memory[92][0] ),
    .I1(\u_cpu.rf_ram.memory[93][0] ),
    .I2(\u_cpu.rf_ram.memory[94][0] ),
    .I3(\u_cpu.rf_ram.memory[95][0] ),
    .S0(_01762_),
    .S1(_01763_),
    .Z(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06148_ (.A1(_01761_),
    .A2(_01764_),
    .ZN(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06149_ (.I(_01671_),
    .Z(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06150_ (.I(_01704_),
    .Z(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06151_ (.I(_01675_),
    .Z(_01768_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06152_ (.I0(\u_cpu.rf_ram.memory[88][0] ),
    .I1(\u_cpu.rf_ram.memory[89][0] ),
    .I2(\u_cpu.rf_ram.memory[90][0] ),
    .I3(\u_cpu.rf_ram.memory[91][0] ),
    .S0(_01767_),
    .S1(_01768_),
    .Z(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06153_ (.I(_01418_),
    .Z(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06154_ (.A1(_01766_),
    .A2(_01769_),
    .B(_01770_),
    .ZN(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06155_ (.I(_01702_),
    .Z(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06156_ (.I(_01685_),
    .Z(_01773_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06157_ (.I(_01652_),
    .Z(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06158_ (.I0(\u_cpu.rf_ram.memory[80][0] ),
    .I1(\u_cpu.rf_ram.memory[81][0] ),
    .I2(\u_cpu.rf_ram.memory[82][0] ),
    .I3(\u_cpu.rf_ram.memory[83][0] ),
    .S0(_01773_),
    .S1(_01774_),
    .Z(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06159_ (.A1(_01772_),
    .A2(_01775_),
    .ZN(_01776_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06160_ (.I(_01397_),
    .Z(_01777_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06161_ (.I(_01777_),
    .Z(_01778_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06162_ (.I(_01572_),
    .Z(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06163_ (.I(_01632_),
    .Z(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06164_ (.I0(\u_cpu.rf_ram.memory[84][0] ),
    .I1(\u_cpu.rf_ram.memory[85][0] ),
    .I2(\u_cpu.rf_ram.memory[86][0] ),
    .I3(\u_cpu.rf_ram.memory[87][0] ),
    .S0(_01779_),
    .S1(_01780_),
    .Z(_01781_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06165_ (.I(_01627_),
    .Z(_01782_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06166_ (.A1(_01778_),
    .A2(_01781_),
    .B(_01782_),
    .ZN(_01783_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06167_ (.I(_01427_),
    .Z(_01784_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06168_ (.A1(_01765_),
    .A2(_01771_),
    .B1(_01776_),
    .B2(_01783_),
    .C(_01784_),
    .ZN(_01785_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06169_ (.I(_01683_),
    .Z(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06170_ (.I(_01612_),
    .Z(_01787_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06171_ (.I(_01575_),
    .Z(_01788_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06172_ (.I0(\u_cpu.rf_ram.memory[64][0] ),
    .I1(\u_cpu.rf_ram.memory[65][0] ),
    .I2(\u_cpu.rf_ram.memory[66][0] ),
    .I3(\u_cpu.rf_ram.memory[67][0] ),
    .S0(_01787_),
    .S1(_01788_),
    .Z(_01789_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06173_ (.A1(_01786_),
    .A2(_01789_),
    .ZN(_01790_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06174_ (.I(_01777_),
    .Z(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06175_ (.I(_01572_),
    .Z(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06176_ (.I(_01632_),
    .Z(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06177_ (.I0(\u_cpu.rf_ram.memory[68][0] ),
    .I1(\u_cpu.rf_ram.memory[69][0] ),
    .I2(\u_cpu.rf_ram.memory[70][0] ),
    .I3(\u_cpu.rf_ram.memory[71][0] ),
    .S0(_01792_),
    .S1(_01793_),
    .Z(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06178_ (.I(_01627_),
    .Z(_01795_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06179_ (.A1(_01791_),
    .A2(_01794_),
    .B(_01795_),
    .ZN(_01796_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06180_ (.I(_01683_),
    .Z(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06181_ (.I(_01612_),
    .Z(_01798_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06182_ (.I(_01584_),
    .Z(_01799_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06183_ (.I0(\u_cpu.rf_ram.memory[72][0] ),
    .I1(\u_cpu.rf_ram.memory[73][0] ),
    .I2(\u_cpu.rf_ram.memory[74][0] ),
    .I3(\u_cpu.rf_ram.memory[75][0] ),
    .S0(_01798_),
    .S1(_01799_),
    .Z(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06184_ (.A1(_01797_),
    .A2(_01800_),
    .ZN(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06185_ (.I(_01777_),
    .Z(_01802_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06186_ (.I(_01706_),
    .Z(_01803_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06187_ (.I0(\u_cpu.rf_ram.memory[76][0] ),
    .I1(\u_cpu.rf_ram.memory[77][0] ),
    .I2(\u_cpu.rf_ram.memory[78][0] ),
    .I3(\u_cpu.rf_ram.memory[79][0] ),
    .S0(_01582_),
    .S1(_01803_),
    .Z(_01804_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06188_ (.I(_01418_),
    .Z(_01805_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06189_ (.A1(_01802_),
    .A2(_01804_),
    .B(_01805_),
    .ZN(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06190_ (.I(_01606_),
    .Z(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06191_ (.A1(_01790_),
    .A2(_01796_),
    .B1(_01801_),
    .B2(_01806_),
    .C(_01807_),
    .ZN(_01808_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06192_ (.A1(_01760_),
    .A2(_01785_),
    .A3(_01808_),
    .ZN(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06193_ (.I(_01404_),
    .Z(_01810_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06194_ (.A1(_01759_),
    .A2(_01809_),
    .B(_01810_),
    .ZN(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06195_ (.I(_01581_),
    .Z(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06196_ (.I(_01812_),
    .Z(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06197_ (.I(_01813_),
    .Z(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06198_ (.I(_01706_),
    .Z(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06199_ (.I(_01815_),
    .Z(_01816_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06200_ (.I0(\u_cpu.rf_ram.memory[136][0] ),
    .I1(\u_cpu.rf_ram.memory[137][0] ),
    .I2(\u_cpu.rf_ram.memory[138][0] ),
    .I3(\u_cpu.rf_ram.memory[139][0] ),
    .S0(_01814_),
    .S1(_01816_),
    .Z(_01817_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06201_ (.A1(_01400_),
    .A2(_01817_),
    .ZN(_01818_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06202_ (.I(_01568_),
    .Z(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06203_ (.I(_01613_),
    .Z(_01820_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06204_ (.I(_01815_),
    .Z(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06205_ (.I0(\u_cpu.rf_ram.memory[140][0] ),
    .I1(\u_cpu.rf_ram.memory[141][0] ),
    .I2(\u_cpu.rf_ram.memory[142][0] ),
    .I3(\u_cpu.rf_ram.memory[143][0] ),
    .S0(_01820_),
    .S1(_01821_),
    .Z(_01822_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06206_ (.I(_01602_),
    .Z(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06207_ (.A1(_01819_),
    .A2(_01822_),
    .B(_01823_),
    .ZN(_01824_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06208_ (.I(_01610_),
    .Z(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06209_ (.I(_01613_),
    .Z(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06210_ (.I(_01788_),
    .Z(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06211_ (.I0(\u_cpu.rf_ram.memory[128][0] ),
    .I1(\u_cpu.rf_ram.memory[129][0] ),
    .I2(\u_cpu.rf_ram.memory[130][0] ),
    .I3(\u_cpu.rf_ram.memory[131][0] ),
    .S0(_01826_),
    .S1(_01827_),
    .Z(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06212_ (.A1(_01825_),
    .A2(_01828_),
    .ZN(_01829_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06213_ (.I(_01568_),
    .Z(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06214_ (.I(_01613_),
    .Z(_01831_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06215_ (.I(_01788_),
    .Z(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06216_ (.I0(\u_cpu.rf_ram.memory[132][0] ),
    .I1(\u_cpu.rf_ram.memory[133][0] ),
    .I2(\u_cpu.rf_ram.memory[134][0] ),
    .I3(\u_cpu.rf_ram.memory[135][0] ),
    .S0(_01831_),
    .S1(_01832_),
    .Z(_01833_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06217_ (.A1(_01830_),
    .A2(_01833_),
    .B(_01419_),
    .ZN(_01834_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06218_ (.I(_01405_),
    .Z(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _06219_ (.A1(_01818_),
    .A2(_01824_),
    .B1(_01829_),
    .B2(_01834_),
    .C(_01835_),
    .ZN(_01836_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06220_ (.A1(_01811_),
    .A2(_01836_),
    .ZN(_01837_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06221_ (.A1(_01564_),
    .A2(_01714_),
    .B(_01837_),
    .ZN(_00000_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06222_ (.I(_01576_),
    .Z(_01838_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06223_ (.I0(\u_cpu.rf_ram.memory[8][1] ),
    .I1(\u_cpu.rf_ram.memory[9][1] ),
    .I2(\u_cpu.rf_ram.memory[10][1] ),
    .I3(\u_cpu.rf_ram.memory[11][1] ),
    .S0(_01574_),
    .S1(_01838_),
    .Z(_01839_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06224_ (.A1(_01570_),
    .A2(_01839_),
    .ZN(_01840_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06225_ (.I(_01584_),
    .Z(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06226_ (.I0(\u_cpu.rf_ram.memory[12][1] ),
    .I1(\u_cpu.rf_ram.memory[13][1] ),
    .I2(\u_cpu.rf_ram.memory[14][1] ),
    .I3(\u_cpu.rf_ram.memory[15][1] ),
    .S0(_01583_),
    .S1(_01841_),
    .Z(_01842_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06227_ (.A1(_01580_),
    .A2(_01842_),
    .B(_01588_),
    .ZN(_01843_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06228_ (.I0(\u_cpu.rf_ram.memory[4][1] ),
    .I1(\u_cpu.rf_ram.memory[5][1] ),
    .I2(\u_cpu.rf_ram.memory[6][1] ),
    .I3(\u_cpu.rf_ram.memory[7][1] ),
    .S0(_01591_),
    .S1(_01592_),
    .Z(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06229_ (.A1(_01590_),
    .A2(_01844_),
    .ZN(_01845_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06230_ (.I0(\u_cpu.rf_ram.memory[0][1] ),
    .I1(\u_cpu.rf_ram.memory[1][1] ),
    .I2(\u_cpu.rf_ram.memory[2][1] ),
    .I3(\u_cpu.rf_ram.memory[3][1] ),
    .S0(_01598_),
    .S1(_01599_),
    .Z(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06231_ (.A1(_01597_),
    .A2(_01846_),
    .B(_01603_),
    .ZN(_01847_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06232_ (.A1(_01840_),
    .A2(_01843_),
    .B1(_01845_),
    .B2(_01847_),
    .C(_01607_),
    .ZN(_01848_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06233_ (.I(_01573_),
    .Z(_01849_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06234_ (.I0(\u_cpu.rf_ram.memory[20][1] ),
    .I1(\u_cpu.rf_ram.memory[21][1] ),
    .I2(\u_cpu.rf_ram.memory[22][1] ),
    .I3(\u_cpu.rf_ram.memory[23][1] ),
    .S0(_01849_),
    .S1(_01616_),
    .Z(_01850_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06235_ (.A1(_01611_),
    .A2(_01850_),
    .ZN(_01851_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06236_ (.I(_01621_),
    .Z(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06237_ (.I0(\u_cpu.rf_ram.memory[16][1] ),
    .I1(\u_cpu.rf_ram.memory[17][1] ),
    .I2(\u_cpu.rf_ram.memory[18][1] ),
    .I3(\u_cpu.rf_ram.memory[19][1] ),
    .S0(_01852_),
    .S1(_01625_),
    .Z(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06238_ (.A1(_01619_),
    .A2(_01853_),
    .B(_01628_),
    .ZN(_01854_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06239_ (.I0(\u_cpu.rf_ram.memory[28][1] ),
    .I1(\u_cpu.rf_ram.memory[29][1] ),
    .I2(\u_cpu.rf_ram.memory[30][1] ),
    .I3(\u_cpu.rf_ram.memory[31][1] ),
    .S0(_01631_),
    .S1(_01634_),
    .Z(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06240_ (.A1(_01630_),
    .A2(_01855_),
    .ZN(_01856_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06241_ (.I(_01596_),
    .Z(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06242_ (.I0(\u_cpu.rf_ram.memory[24][1] ),
    .I1(\u_cpu.rf_ram.memory[25][1] ),
    .I2(\u_cpu.rf_ram.memory[26][1] ),
    .I3(\u_cpu.rf_ram.memory[27][1] ),
    .S0(_01640_),
    .S1(_01642_),
    .Z(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06243_ (.I(_01587_),
    .Z(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06244_ (.A1(_01857_),
    .A2(_01858_),
    .B(_01859_),
    .ZN(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06245_ (.A1(_01851_),
    .A2(_01854_),
    .B1(_01856_),
    .B2(_01860_),
    .C(_01428_),
    .ZN(_01861_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06246_ (.I(_01422_),
    .Z(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06247_ (.I(_01650_),
    .Z(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06248_ (.I0(\u_cpu.rf_ram.memory[52][1] ),
    .I1(\u_cpu.rf_ram.memory[53][1] ),
    .I2(\u_cpu.rf_ram.memory[54][1] ),
    .I3(\u_cpu.rf_ram.memory[55][1] ),
    .S0(_01863_),
    .S1(_01653_),
    .Z(_01864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06249_ (.A1(_01649_),
    .A2(_01864_),
    .ZN(_01865_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06250_ (.I0(\u_cpu.rf_ram.memory[48][1] ),
    .I1(\u_cpu.rf_ram.memory[49][1] ),
    .I2(\u_cpu.rf_ram.memory[50][1] ),
    .I3(\u_cpu.rf_ram.memory[51][1] ),
    .S0(_01657_),
    .S1(_01660_),
    .Z(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06251_ (.I(_01601_),
    .Z(_01867_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06252_ (.A1(_01656_),
    .A2(_01866_),
    .B(_01867_),
    .ZN(_01868_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06253_ (.I0(\u_cpu.rf_ram.memory[60][1] ),
    .I1(\u_cpu.rf_ram.memory[61][1] ),
    .I2(\u_cpu.rf_ram.memory[62][1] ),
    .I3(\u_cpu.rf_ram.memory[63][1] ),
    .S0(_01639_),
    .S1(_01668_),
    .Z(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06254_ (.A1(_01666_),
    .A2(_01869_),
    .ZN(_01870_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06255_ (.I(_01673_),
    .Z(_01871_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06256_ (.I0(\u_cpu.rf_ram.memory[56][1] ),
    .I1(\u_cpu.rf_ram.memory[57][1] ),
    .I2(\u_cpu.rf_ram.memory[58][1] ),
    .I3(\u_cpu.rf_ram.memory[59][1] ),
    .S0(_01871_),
    .S1(_01676_),
    .Z(_01872_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06257_ (.I(_01678_),
    .Z(_01873_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06258_ (.A1(_01672_),
    .A2(_01872_),
    .B(_01873_),
    .ZN(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06259_ (.A1(_01865_),
    .A2(_01868_),
    .B1(_01870_),
    .B2(_01874_),
    .C(_01681_),
    .ZN(_01875_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06260_ (.I(_01683_),
    .Z(_01876_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06261_ (.I0(\u_cpu.rf_ram.memory[40][1] ),
    .I1(\u_cpu.rf_ram.memory[41][1] ),
    .I2(\u_cpu.rf_ram.memory[42][1] ),
    .I3(\u_cpu.rf_ram.memory[43][1] ),
    .S0(_01686_),
    .S1(_01688_),
    .Z(_01877_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06262_ (.A1(_01876_),
    .A2(_01877_),
    .ZN(_01878_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06263_ (.I(_01659_),
    .Z(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06264_ (.I0(\u_cpu.rf_ram.memory[44][1] ),
    .I1(\u_cpu.rf_ram.memory[45][1] ),
    .I2(\u_cpu.rf_ram.memory[46][1] ),
    .I3(\u_cpu.rf_ram.memory[47][1] ),
    .S0(_01692_),
    .S1(_01879_),
    .Z(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06265_ (.A1(_01691_),
    .A2(_01880_),
    .B(_01695_),
    .ZN(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06266_ (.I(_01665_),
    .Z(_01882_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06267_ (.I0(\u_cpu.rf_ram.memory[36][1] ),
    .I1(\u_cpu.rf_ram.memory[37][1] ),
    .I2(\u_cpu.rf_ram.memory[38][1] ),
    .I3(\u_cpu.rf_ram.memory[39][1] ),
    .S0(_01698_),
    .S1(_01699_),
    .Z(_01883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06268_ (.A1(_01882_),
    .A2(_01883_),
    .ZN(_01884_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06269_ (.I0(\u_cpu.rf_ram.memory[32][1] ),
    .I1(\u_cpu.rf_ram.memory[33][1] ),
    .I2(\u_cpu.rf_ram.memory[34][1] ),
    .I3(\u_cpu.rf_ram.memory[35][1] ),
    .S0(_01705_),
    .S1(_01707_),
    .Z(_01885_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06270_ (.A1(_01703_),
    .A2(_01885_),
    .B(_01709_),
    .ZN(_01886_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06271_ (.A1(_01878_),
    .A2(_01881_),
    .B1(_01884_),
    .B2(_01886_),
    .C(_01711_),
    .ZN(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06272_ (.A1(_01862_),
    .A2(_01875_),
    .A3(_01887_),
    .Z(_01888_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06273_ (.A1(_01566_),
    .A2(_01848_),
    .A3(_01861_),
    .B(_01888_),
    .ZN(_01889_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06274_ (.I0(\u_cpu.rf_ram.memory[108][1] ),
    .I1(\u_cpu.rf_ram.memory[109][1] ),
    .I2(\u_cpu.rf_ram.memory[110][1] ),
    .I3(\u_cpu.rf_ram.memory[111][1] ),
    .S0(_01716_),
    .S1(_01717_),
    .Z(_01890_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06275_ (.A1(_01715_),
    .A2(_01890_),
    .ZN(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06276_ (.I(_01659_),
    .Z(_01892_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06277_ (.I0(\u_cpu.rf_ram.memory[104][1] ),
    .I1(\u_cpu.rf_ram.memory[105][1] ),
    .I2(\u_cpu.rf_ram.memory[106][1] ),
    .I3(\u_cpu.rf_ram.memory[107][1] ),
    .S0(_01721_),
    .S1(_01892_),
    .Z(_01893_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06278_ (.A1(_01720_),
    .A2(_01893_),
    .B(_01723_),
    .ZN(_01894_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06279_ (.I(_01667_),
    .Z(_01895_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06280_ (.I0(\u_cpu.rf_ram.memory[100][1] ),
    .I1(\u_cpu.rf_ram.memory[101][1] ),
    .I2(\u_cpu.rf_ram.memory[102][1] ),
    .I3(\u_cpu.rf_ram.memory[103][1] ),
    .S0(_01621_),
    .S1(_01895_),
    .Z(_01896_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06281_ (.A1(_01725_),
    .A2(_01896_),
    .ZN(_01897_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06282_ (.I0(\u_cpu.rf_ram.memory[96][1] ),
    .I1(\u_cpu.rf_ram.memory[97][1] ),
    .I2(\u_cpu.rf_ram.memory[98][1] ),
    .I3(\u_cpu.rf_ram.memory[99][1] ),
    .S0(_01729_),
    .S1(_01641_),
    .Z(_01898_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06283_ (.A1(_01728_),
    .A2(_01898_),
    .B(_01731_),
    .ZN(_01899_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06284_ (.I(_01605_),
    .Z(_01900_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06285_ (.A1(_01891_),
    .A2(_01894_),
    .B1(_01897_),
    .B2(_01899_),
    .C(_01900_),
    .ZN(_01901_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06286_ (.I0(\u_cpu.rf_ram.memory[124][1] ),
    .I1(\u_cpu.rf_ram.memory[125][1] ),
    .I2(\u_cpu.rf_ram.memory[126][1] ),
    .I3(\u_cpu.rf_ram.memory[127][1] ),
    .S0(_01736_),
    .S1(_01737_),
    .Z(_01902_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06287_ (.A1(_01735_),
    .A2(_01902_),
    .ZN(_01903_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06288_ (.I(_01671_),
    .Z(_01904_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06289_ (.I(_01675_),
    .Z(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06290_ (.I0(\u_cpu.rf_ram.memory[120][1] ),
    .I1(\u_cpu.rf_ram.memory[121][1] ),
    .I2(\u_cpu.rf_ram.memory[122][1] ),
    .I3(\u_cpu.rf_ram.memory[123][1] ),
    .S0(_01741_),
    .S1(_01905_),
    .Z(_01906_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06291_ (.A1(_01904_),
    .A2(_01906_),
    .B(_01744_),
    .ZN(_01907_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06292_ (.I(_01652_),
    .Z(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06293_ (.I0(\u_cpu.rf_ram.memory[112][1] ),
    .I1(\u_cpu.rf_ram.memory[113][1] ),
    .I2(\u_cpu.rf_ram.memory[114][1] ),
    .I3(\u_cpu.rf_ram.memory[115][1] ),
    .S0(_01747_),
    .S1(_01908_),
    .Z(_01909_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06294_ (.A1(_01746_),
    .A2(_01909_),
    .ZN(_01910_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06295_ (.I0(\u_cpu.rf_ram.memory[116][1] ),
    .I1(\u_cpu.rf_ram.memory[117][1] ),
    .I2(\u_cpu.rf_ram.memory[118][1] ),
    .I3(\u_cpu.rf_ram.memory[119][1] ),
    .S0(_01752_),
    .S1(_01753_),
    .Z(_01911_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06296_ (.A1(_01751_),
    .A2(_01911_),
    .B(_01755_),
    .ZN(_01912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06297_ (.A1(_01903_),
    .A2(_01907_),
    .B1(_01910_),
    .B2(_01912_),
    .C(_01757_),
    .ZN(_01913_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06298_ (.A1(_01423_),
    .A2(_01901_),
    .A3(_01913_),
    .ZN(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06299_ (.I(_01687_),
    .Z(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06300_ (.I0(\u_cpu.rf_ram.memory[92][1] ),
    .I1(\u_cpu.rf_ram.memory[93][1] ),
    .I2(\u_cpu.rf_ram.memory[94][1] ),
    .I3(\u_cpu.rf_ram.memory[95][1] ),
    .S0(_01762_),
    .S1(_01915_),
    .Z(_01916_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06301_ (.A1(_01761_),
    .A2(_01916_),
    .ZN(_01917_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06302_ (.I0(\u_cpu.rf_ram.memory[88][1] ),
    .I1(\u_cpu.rf_ram.memory[89][1] ),
    .I2(\u_cpu.rf_ram.memory[90][1] ),
    .I3(\u_cpu.rf_ram.memory[91][1] ),
    .S0(_01767_),
    .S1(_01768_),
    .Z(_01918_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06303_ (.A1(_01766_),
    .A2(_01918_),
    .B(_01770_),
    .ZN(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06304_ (.I0(\u_cpu.rf_ram.memory[80][1] ),
    .I1(\u_cpu.rf_ram.memory[81][1] ),
    .I2(\u_cpu.rf_ram.memory[82][1] ),
    .I3(\u_cpu.rf_ram.memory[83][1] ),
    .S0(_01773_),
    .S1(_01774_),
    .Z(_01920_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06305_ (.A1(_01772_),
    .A2(_01920_),
    .ZN(_01921_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06306_ (.I(_01572_),
    .Z(_01922_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06307_ (.I0(\u_cpu.rf_ram.memory[84][1] ),
    .I1(\u_cpu.rf_ram.memory[85][1] ),
    .I2(\u_cpu.rf_ram.memory[86][1] ),
    .I3(\u_cpu.rf_ram.memory[87][1] ),
    .S0(_01922_),
    .S1(_01780_),
    .Z(_01923_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06308_ (.A1(_01778_),
    .A2(_01923_),
    .B(_01782_),
    .ZN(_01924_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06309_ (.I(_01426_),
    .Z(_01925_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06310_ (.A1(_01917_),
    .A2(_01919_),
    .B1(_01921_),
    .B2(_01924_),
    .C(_01925_),
    .ZN(_01926_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06311_ (.I0(\u_cpu.rf_ram.memory[64][1] ),
    .I1(\u_cpu.rf_ram.memory[65][1] ),
    .I2(\u_cpu.rf_ram.memory[66][1] ),
    .I3(\u_cpu.rf_ram.memory[67][1] ),
    .S0(_01787_),
    .S1(_01788_),
    .Z(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06312_ (.A1(_01786_),
    .A2(_01927_),
    .ZN(_01928_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06313_ (.I(_01777_),
    .Z(_01929_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06314_ (.I(_01632_),
    .Z(_01930_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06315_ (.I0(\u_cpu.rf_ram.memory[68][1] ),
    .I1(\u_cpu.rf_ram.memory[69][1] ),
    .I2(\u_cpu.rf_ram.memory[70][1] ),
    .I3(\u_cpu.rf_ram.memory[71][1] ),
    .S0(_01792_),
    .S1(_01930_),
    .Z(_01931_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06316_ (.I(_01627_),
    .Z(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06317_ (.A1(_01929_),
    .A2(_01931_),
    .B(_01932_),
    .ZN(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06318_ (.I(_01612_),
    .Z(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06319_ (.I0(\u_cpu.rf_ram.memory[72][1] ),
    .I1(\u_cpu.rf_ram.memory[73][1] ),
    .I2(\u_cpu.rf_ram.memory[74][1] ),
    .I3(\u_cpu.rf_ram.memory[75][1] ),
    .S0(_01934_),
    .S1(_01799_),
    .Z(_01935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06320_ (.A1(_01797_),
    .A2(_01935_),
    .ZN(_01936_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06321_ (.I0(\u_cpu.rf_ram.memory[76][1] ),
    .I1(\u_cpu.rf_ram.memory[77][1] ),
    .I2(\u_cpu.rf_ram.memory[78][1] ),
    .I3(\u_cpu.rf_ram.memory[79][1] ),
    .S0(_01582_),
    .S1(_01803_),
    .Z(_01937_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06322_ (.A1(_01802_),
    .A2(_01937_),
    .B(_01805_),
    .ZN(_01938_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06323_ (.A1(_01928_),
    .A2(_01933_),
    .B1(_01936_),
    .B2(_01938_),
    .C(_01807_),
    .ZN(_01939_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06324_ (.A1(_01760_),
    .A2(_01926_),
    .A3(_01939_),
    .ZN(_01940_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06325_ (.A1(_01914_),
    .A2(_01940_),
    .B(_01810_),
    .ZN(_01941_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06326_ (.I(_01815_),
    .Z(_01942_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06327_ (.I0(\u_cpu.rf_ram.memory[136][1] ),
    .I1(\u_cpu.rf_ram.memory[137][1] ),
    .I2(\u_cpu.rf_ram.memory[138][1] ),
    .I3(\u_cpu.rf_ram.memory[139][1] ),
    .S0(_01814_),
    .S1(_01942_),
    .Z(_01943_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06328_ (.A1(_01400_),
    .A2(_01943_),
    .ZN(_01944_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06329_ (.I0(\u_cpu.rf_ram.memory[140][1] ),
    .I1(\u_cpu.rf_ram.memory[141][1] ),
    .I2(\u_cpu.rf_ram.memory[142][1] ),
    .I3(\u_cpu.rf_ram.memory[143][1] ),
    .S0(_01820_),
    .S1(_01821_),
    .Z(_01945_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06330_ (.A1(_01819_),
    .A2(_01945_),
    .B(_01823_),
    .ZN(_01946_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06331_ (.I(_01610_),
    .Z(_01947_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06332_ (.I0(\u_cpu.rf_ram.memory[128][1] ),
    .I1(\u_cpu.rf_ram.memory[129][1] ),
    .I2(\u_cpu.rf_ram.memory[130][1] ),
    .I3(\u_cpu.rf_ram.memory[131][1] ),
    .S0(_01826_),
    .S1(_01827_),
    .Z(_01948_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06333_ (.A1(_01947_),
    .A2(_01948_),
    .ZN(_01949_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06334_ (.I0(\u_cpu.rf_ram.memory[132][1] ),
    .I1(\u_cpu.rf_ram.memory[133][1] ),
    .I2(\u_cpu.rf_ram.memory[134][1] ),
    .I3(\u_cpu.rf_ram.memory[135][1] ),
    .S0(_01831_),
    .S1(_01832_),
    .Z(_01950_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06335_ (.A1(_01830_),
    .A2(_01950_),
    .B(_01419_),
    .ZN(_01951_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _06336_ (.A1(_01944_),
    .A2(_01946_),
    .B1(_01949_),
    .B2(_01951_),
    .C(_01835_),
    .ZN(_01952_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06337_ (.A1(_01941_),
    .A2(_01952_),
    .ZN(_01953_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06338_ (.A1(_01564_),
    .A2(_01889_),
    .B(_01953_),
    .ZN(_00001_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06339_ (.I0(\u_cpu.rf_ram.memory[8][2] ),
    .I1(\u_cpu.rf_ram.memory[9][2] ),
    .I2(\u_cpu.rf_ram.memory[10][2] ),
    .I3(\u_cpu.rf_ram.memory[11][2] ),
    .S0(_01574_),
    .S1(_01838_),
    .Z(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06340_ (.A1(_01570_),
    .A2(_01954_),
    .ZN(_01955_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06341_ (.I0(\u_cpu.rf_ram.memory[12][2] ),
    .I1(\u_cpu.rf_ram.memory[13][2] ),
    .I2(\u_cpu.rf_ram.memory[14][2] ),
    .I3(\u_cpu.rf_ram.memory[15][2] ),
    .S0(_01583_),
    .S1(_01841_),
    .Z(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06342_ (.A1(_01580_),
    .A2(_01956_),
    .B(_01588_),
    .ZN(_01957_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06343_ (.I(_01398_),
    .Z(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06344_ (.I(_01787_),
    .Z(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06345_ (.I0(\u_cpu.rf_ram.memory[4][2] ),
    .I1(\u_cpu.rf_ram.memory[5][2] ),
    .I2(\u_cpu.rf_ram.memory[6][2] ),
    .I3(\u_cpu.rf_ram.memory[7][2] ),
    .S0(_01959_),
    .S1(_01592_),
    .Z(_01960_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06346_ (.A1(_01958_),
    .A2(_01960_),
    .ZN(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06347_ (.I0(\u_cpu.rf_ram.memory[0][2] ),
    .I1(\u_cpu.rf_ram.memory[1][2] ),
    .I2(\u_cpu.rf_ram.memory[2][2] ),
    .I3(\u_cpu.rf_ram.memory[3][2] ),
    .S0(_01598_),
    .S1(_01599_),
    .Z(_01962_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06348_ (.A1(_01597_),
    .A2(_01962_),
    .B(_01603_),
    .ZN(_01963_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06349_ (.A1(_01955_),
    .A2(_01957_),
    .B1(_01961_),
    .B2(_01963_),
    .C(_01607_),
    .ZN(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06350_ (.I(_01615_),
    .Z(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06351_ (.I0(\u_cpu.rf_ram.memory[20][2] ),
    .I1(\u_cpu.rf_ram.memory[21][2] ),
    .I2(\u_cpu.rf_ram.memory[22][2] ),
    .I3(\u_cpu.rf_ram.memory[23][2] ),
    .S0(_01849_),
    .S1(_01965_),
    .Z(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06352_ (.A1(_01611_),
    .A2(_01966_),
    .ZN(_01967_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06353_ (.I(_01624_),
    .Z(_01968_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06354_ (.I0(\u_cpu.rf_ram.memory[16][2] ),
    .I1(\u_cpu.rf_ram.memory[17][2] ),
    .I2(\u_cpu.rf_ram.memory[18][2] ),
    .I3(\u_cpu.rf_ram.memory[19][2] ),
    .S0(_01852_),
    .S1(_01968_),
    .Z(_01969_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06355_ (.I(_01602_),
    .Z(_01970_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06356_ (.A1(_01619_),
    .A2(_01969_),
    .B(_01970_),
    .ZN(_01971_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06357_ (.I0(\u_cpu.rf_ram.memory[28][2] ),
    .I1(\u_cpu.rf_ram.memory[29][2] ),
    .I2(\u_cpu.rf_ram.memory[30][2] ),
    .I3(\u_cpu.rf_ram.memory[31][2] ),
    .S0(_01631_),
    .S1(_01634_),
    .Z(_01972_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06358_ (.A1(_01630_),
    .A2(_01972_),
    .ZN(_01973_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06359_ (.I0(\u_cpu.rf_ram.memory[24][2] ),
    .I1(\u_cpu.rf_ram.memory[25][2] ),
    .I2(\u_cpu.rf_ram.memory[26][2] ),
    .I3(\u_cpu.rf_ram.memory[27][2] ),
    .S0(_01640_),
    .S1(_01642_),
    .Z(_01974_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06360_ (.A1(_01857_),
    .A2(_01974_),
    .B(_01859_),
    .ZN(_01975_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06361_ (.A1(_01967_),
    .A2(_01971_),
    .B1(_01973_),
    .B2(_01975_),
    .C(_01428_),
    .ZN(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06362_ (.I0(\u_cpu.rf_ram.memory[52][2] ),
    .I1(\u_cpu.rf_ram.memory[53][2] ),
    .I2(\u_cpu.rf_ram.memory[54][2] ),
    .I3(\u_cpu.rf_ram.memory[55][2] ),
    .S0(_01863_),
    .S1(_01653_),
    .Z(_01977_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06363_ (.A1(_01649_),
    .A2(_01977_),
    .ZN(_01978_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06364_ (.I0(\u_cpu.rf_ram.memory[48][2] ),
    .I1(\u_cpu.rf_ram.memory[49][2] ),
    .I2(\u_cpu.rf_ram.memory[50][2] ),
    .I3(\u_cpu.rf_ram.memory[51][2] ),
    .S0(_01657_),
    .S1(_01660_),
    .Z(_01979_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06365_ (.A1(_01656_),
    .A2(_01979_),
    .B(_01867_),
    .ZN(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06366_ (.I0(\u_cpu.rf_ram.memory[60][2] ),
    .I1(\u_cpu.rf_ram.memory[61][2] ),
    .I2(\u_cpu.rf_ram.memory[62][2] ),
    .I3(\u_cpu.rf_ram.memory[63][2] ),
    .S0(_01639_),
    .S1(_01668_),
    .Z(_01981_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06367_ (.A1(_01666_),
    .A2(_01981_),
    .ZN(_01982_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06368_ (.I0(\u_cpu.rf_ram.memory[56][2] ),
    .I1(\u_cpu.rf_ram.memory[57][2] ),
    .I2(\u_cpu.rf_ram.memory[58][2] ),
    .I3(\u_cpu.rf_ram.memory[59][2] ),
    .S0(_01871_),
    .S1(_01676_),
    .Z(_01983_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06369_ (.A1(_01672_),
    .A2(_01983_),
    .B(_01873_),
    .ZN(_01984_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06370_ (.A1(_01978_),
    .A2(_01980_),
    .B1(_01982_),
    .B2(_01984_),
    .C(_01681_),
    .ZN(_01985_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06371_ (.I0(\u_cpu.rf_ram.memory[40][2] ),
    .I1(\u_cpu.rf_ram.memory[41][2] ),
    .I2(\u_cpu.rf_ram.memory[42][2] ),
    .I3(\u_cpu.rf_ram.memory[43][2] ),
    .S0(_01686_),
    .S1(_01688_),
    .Z(_01986_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06372_ (.A1(_01876_),
    .A2(_01986_),
    .ZN(_01987_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06373_ (.I(_01609_),
    .Z(_01988_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06374_ (.I0(\u_cpu.rf_ram.memory[44][2] ),
    .I1(\u_cpu.rf_ram.memory[45][2] ),
    .I2(\u_cpu.rf_ram.memory[46][2] ),
    .I3(\u_cpu.rf_ram.memory[47][2] ),
    .S0(_01692_),
    .S1(_01879_),
    .Z(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06375_ (.A1(_01988_),
    .A2(_01989_),
    .B(_01695_),
    .ZN(_01990_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06376_ (.I0(\u_cpu.rf_ram.memory[36][2] ),
    .I1(\u_cpu.rf_ram.memory[37][2] ),
    .I2(\u_cpu.rf_ram.memory[38][2] ),
    .I3(\u_cpu.rf_ram.memory[39][2] ),
    .S0(_01698_),
    .S1(_01699_),
    .Z(_01991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06377_ (.A1(_01882_),
    .A2(_01991_),
    .ZN(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06378_ (.I(_01702_),
    .Z(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06379_ (.I(_01706_),
    .Z(_01994_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06380_ (.I0(\u_cpu.rf_ram.memory[32][2] ),
    .I1(\u_cpu.rf_ram.memory[33][2] ),
    .I2(\u_cpu.rf_ram.memory[34][2] ),
    .I3(\u_cpu.rf_ram.memory[35][2] ),
    .S0(_01705_),
    .S1(_01994_),
    .Z(_01995_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06381_ (.I(_01662_),
    .Z(_01996_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06382_ (.A1(_01993_),
    .A2(_01995_),
    .B(_01996_),
    .ZN(_01997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06383_ (.A1(_01987_),
    .A2(_01990_),
    .B1(_01992_),
    .B2(_01997_),
    .C(_01711_),
    .ZN(_01998_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06384_ (.A1(_01862_),
    .A2(_01985_),
    .A3(_01998_),
    .Z(_01999_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06385_ (.A1(_01566_),
    .A2(_01964_),
    .A3(_01976_),
    .B(_01999_),
    .ZN(_02000_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06386_ (.I(_01638_),
    .Z(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06387_ (.I0(\u_cpu.rf_ram.memory[108][2] ),
    .I1(\u_cpu.rf_ram.memory[109][2] ),
    .I2(\u_cpu.rf_ram.memory[110][2] ),
    .I3(\u_cpu.rf_ram.memory[111][2] ),
    .S0(_02001_),
    .S1(_01717_),
    .Z(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06388_ (.A1(_01715_),
    .A2(_02002_),
    .ZN(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06389_ (.I(_01595_),
    .Z(_02004_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06390_ (.I(_01620_),
    .Z(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06391_ (.I0(\u_cpu.rf_ram.memory[104][2] ),
    .I1(\u_cpu.rf_ram.memory[105][2] ),
    .I2(\u_cpu.rf_ram.memory[106][2] ),
    .I3(\u_cpu.rf_ram.memory[107][2] ),
    .S0(_02005_),
    .S1(_01892_),
    .Z(_02006_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06392_ (.A1(_02004_),
    .A2(_02006_),
    .B(_01723_),
    .ZN(_02007_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06393_ (.I(_01777_),
    .Z(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06394_ (.I0(\u_cpu.rf_ram.memory[100][2] ),
    .I1(\u_cpu.rf_ram.memory[101][2] ),
    .I2(\u_cpu.rf_ram.memory[102][2] ),
    .I3(\u_cpu.rf_ram.memory[103][2] ),
    .S0(_01621_),
    .S1(_01895_),
    .Z(_02009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06395_ (.A1(_02008_),
    .A2(_02009_),
    .ZN(_02010_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06396_ (.I0(\u_cpu.rf_ram.memory[96][2] ),
    .I1(\u_cpu.rf_ram.memory[97][2] ),
    .I2(\u_cpu.rf_ram.memory[98][2] ),
    .I3(\u_cpu.rf_ram.memory[99][2] ),
    .S0(_01729_),
    .S1(_01641_),
    .Z(_02011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06397_ (.A1(_01728_),
    .A2(_02011_),
    .B(_01731_),
    .ZN(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06398_ (.A1(_02003_),
    .A2(_02007_),
    .B1(_02010_),
    .B2(_02012_),
    .C(_01900_),
    .ZN(_02013_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06399_ (.I(_01648_),
    .Z(_02014_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06400_ (.I(_01685_),
    .Z(_02015_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06401_ (.I0(\u_cpu.rf_ram.memory[124][2] ),
    .I1(\u_cpu.rf_ram.memory[125][2] ),
    .I2(\u_cpu.rf_ram.memory[126][2] ),
    .I3(\u_cpu.rf_ram.memory[127][2] ),
    .S0(_02015_),
    .S1(_01737_),
    .Z(_02016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06402_ (.A1(_02014_),
    .A2(_02016_),
    .ZN(_02017_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06403_ (.I0(\u_cpu.rf_ram.memory[120][2] ),
    .I1(\u_cpu.rf_ram.memory[121][2] ),
    .I2(\u_cpu.rf_ram.memory[122][2] ),
    .I3(\u_cpu.rf_ram.memory[123][2] ),
    .S0(_01741_),
    .S1(_01905_),
    .Z(_02018_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06404_ (.A1(_01904_),
    .A2(_02018_),
    .B(_01744_),
    .ZN(_02019_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06405_ (.I0(\u_cpu.rf_ram.memory[112][2] ),
    .I1(\u_cpu.rf_ram.memory[113][2] ),
    .I2(\u_cpu.rf_ram.memory[114][2] ),
    .I3(\u_cpu.rf_ram.memory[115][2] ),
    .S0(_01747_),
    .S1(_01908_),
    .Z(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06406_ (.A1(_01746_),
    .A2(_02020_),
    .ZN(_02021_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06407_ (.I0(\u_cpu.rf_ram.memory[116][2] ),
    .I1(\u_cpu.rf_ram.memory[117][2] ),
    .I2(\u_cpu.rf_ram.memory[118][2] ),
    .I3(\u_cpu.rf_ram.memory[119][2] ),
    .S0(_01752_),
    .S1(_01753_),
    .Z(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06408_ (.A1(_01751_),
    .A2(_02022_),
    .B(_01755_),
    .ZN(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06409_ (.A1(_02017_),
    .A2(_02019_),
    .B1(_02021_),
    .B2(_02023_),
    .C(_01757_),
    .ZN(_02024_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06410_ (.A1(_01423_),
    .A2(_02013_),
    .A3(_02024_),
    .ZN(_02025_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06411_ (.I(_01565_),
    .Z(_02026_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06412_ (.I0(\u_cpu.rf_ram.memory[92][2] ),
    .I1(\u_cpu.rf_ram.memory[93][2] ),
    .I2(\u_cpu.rf_ram.memory[94][2] ),
    .I3(\u_cpu.rf_ram.memory[95][2] ),
    .S0(_01762_),
    .S1(_01915_),
    .Z(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06413_ (.A1(_01761_),
    .A2(_02027_),
    .ZN(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06414_ (.I(_01704_),
    .Z(_02029_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06415_ (.I0(\u_cpu.rf_ram.memory[88][2] ),
    .I1(\u_cpu.rf_ram.memory[89][2] ),
    .I2(\u_cpu.rf_ram.memory[90][2] ),
    .I3(\u_cpu.rf_ram.memory[91][2] ),
    .S0(_02029_),
    .S1(_01768_),
    .Z(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06416_ (.I(_01678_),
    .Z(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06417_ (.A1(_01766_),
    .A2(_02030_),
    .B(_02031_),
    .ZN(_02032_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06418_ (.I(_01652_),
    .Z(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06419_ (.I0(\u_cpu.rf_ram.memory[80][2] ),
    .I1(\u_cpu.rf_ram.memory[81][2] ),
    .I2(\u_cpu.rf_ram.memory[82][2] ),
    .I3(\u_cpu.rf_ram.memory[83][2] ),
    .S0(_01773_),
    .S1(_02033_),
    .Z(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06420_ (.A1(_01772_),
    .A2(_02034_),
    .ZN(_02035_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06421_ (.I0(\u_cpu.rf_ram.memory[84][2] ),
    .I1(\u_cpu.rf_ram.memory[85][2] ),
    .I2(\u_cpu.rf_ram.memory[86][2] ),
    .I3(\u_cpu.rf_ram.memory[87][2] ),
    .S0(_01922_),
    .S1(_01780_),
    .Z(_02036_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06422_ (.A1(_01778_),
    .A2(_02036_),
    .B(_01782_),
    .ZN(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06423_ (.A1(_02028_),
    .A2(_02032_),
    .B1(_02035_),
    .B2(_02037_),
    .C(_01925_),
    .ZN(_02038_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06424_ (.I(_01683_),
    .Z(_02039_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06425_ (.I(_01584_),
    .Z(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06426_ (.I0(\u_cpu.rf_ram.memory[64][2] ),
    .I1(\u_cpu.rf_ram.memory[65][2] ),
    .I2(\u_cpu.rf_ram.memory[66][2] ),
    .I3(\u_cpu.rf_ram.memory[67][2] ),
    .S0(_01787_),
    .S1(_02040_),
    .Z(_02041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06427_ (.A1(_02039_),
    .A2(_02041_),
    .ZN(_02042_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06428_ (.I0(\u_cpu.rf_ram.memory[68][2] ),
    .I1(\u_cpu.rf_ram.memory[69][2] ),
    .I2(\u_cpu.rf_ram.memory[70][2] ),
    .I3(\u_cpu.rf_ram.memory[71][2] ),
    .S0(_01792_),
    .S1(_01930_),
    .Z(_02043_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06429_ (.A1(_01929_),
    .A2(_02043_),
    .B(_01932_),
    .ZN(_02044_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06430_ (.I0(\u_cpu.rf_ram.memory[72][2] ),
    .I1(\u_cpu.rf_ram.memory[73][2] ),
    .I2(\u_cpu.rf_ram.memory[74][2] ),
    .I3(\u_cpu.rf_ram.memory[75][2] ),
    .S0(_01934_),
    .S1(_01799_),
    .Z(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06431_ (.A1(_01797_),
    .A2(_02045_),
    .ZN(_02046_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06432_ (.I(_01572_),
    .Z(_02047_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06433_ (.I0(\u_cpu.rf_ram.memory[76][2] ),
    .I1(\u_cpu.rf_ram.memory[77][2] ),
    .I2(\u_cpu.rf_ram.memory[78][2] ),
    .I3(\u_cpu.rf_ram.memory[79][2] ),
    .S0(_02047_),
    .S1(_01803_),
    .Z(_02048_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06434_ (.A1(_01802_),
    .A2(_02048_),
    .B(_01805_),
    .ZN(_02049_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06435_ (.I(_01606_),
    .Z(_02050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06436_ (.A1(_02042_),
    .A2(_02044_),
    .B1(_02046_),
    .B2(_02049_),
    .C(_02050_),
    .ZN(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06437_ (.A1(_02026_),
    .A2(_02038_),
    .A3(_02051_),
    .ZN(_02052_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06438_ (.A1(_02025_),
    .A2(_02052_),
    .B(_01810_),
    .ZN(_02053_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06439_ (.I0(\u_cpu.rf_ram.memory[136][2] ),
    .I1(\u_cpu.rf_ram.memory[137][2] ),
    .I2(\u_cpu.rf_ram.memory[138][2] ),
    .I3(\u_cpu.rf_ram.memory[139][2] ),
    .S0(_01814_),
    .S1(_01942_),
    .Z(_02054_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06440_ (.A1(_01400_),
    .A2(_02054_),
    .ZN(_02055_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06441_ (.I0(\u_cpu.rf_ram.memory[140][2] ),
    .I1(\u_cpu.rf_ram.memory[141][2] ),
    .I2(\u_cpu.rf_ram.memory[142][2] ),
    .I3(\u_cpu.rf_ram.memory[143][2] ),
    .S0(_01820_),
    .S1(_01821_),
    .Z(_02056_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06442_ (.A1(_01819_),
    .A2(_02056_),
    .B(_01823_),
    .ZN(_02057_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06443_ (.I0(\u_cpu.rf_ram.memory[128][2] ),
    .I1(\u_cpu.rf_ram.memory[129][2] ),
    .I2(\u_cpu.rf_ram.memory[130][2] ),
    .I3(\u_cpu.rf_ram.memory[131][2] ),
    .S0(_01826_),
    .S1(_01827_),
    .Z(_02058_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06444_ (.A1(_01947_),
    .A2(_02058_),
    .ZN(_02059_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06445_ (.I(_01568_),
    .Z(_02060_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06446_ (.I(_01613_),
    .Z(_02061_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06447_ (.I0(\u_cpu.rf_ram.memory[132][2] ),
    .I1(\u_cpu.rf_ram.memory[133][2] ),
    .I2(\u_cpu.rf_ram.memory[134][2] ),
    .I3(\u_cpu.rf_ram.memory[135][2] ),
    .S0(_02061_),
    .S1(_01832_),
    .Z(_02062_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06448_ (.A1(_02060_),
    .A2(_02062_),
    .B(_01419_),
    .ZN(_02063_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _06449_ (.A1(_02055_),
    .A2(_02057_),
    .B1(_02059_),
    .B2(_02063_),
    .C(_01835_),
    .ZN(_02064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06450_ (.A1(_02053_),
    .A2(_02064_),
    .ZN(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06451_ (.A1(_01564_),
    .A2(_02000_),
    .B(_02065_),
    .ZN(_00002_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06452_ (.I0(\u_cpu.rf_ram.memory[8][3] ),
    .I1(\u_cpu.rf_ram.memory[9][3] ),
    .I2(\u_cpu.rf_ram.memory[10][3] ),
    .I3(\u_cpu.rf_ram.memory[11][3] ),
    .S0(_01574_),
    .S1(_01838_),
    .Z(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06453_ (.A1(_01570_),
    .A2(_02066_),
    .ZN(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06454_ (.I0(\u_cpu.rf_ram.memory[12][3] ),
    .I1(\u_cpu.rf_ram.memory[13][3] ),
    .I2(\u_cpu.rf_ram.memory[14][3] ),
    .I3(\u_cpu.rf_ram.memory[15][3] ),
    .S0(_01583_),
    .S1(_01841_),
    .Z(_02068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06455_ (.I(_01418_),
    .Z(_02069_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06456_ (.A1(_01580_),
    .A2(_02068_),
    .B(_02069_),
    .ZN(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06457_ (.I(_01803_),
    .Z(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06458_ (.I0(\u_cpu.rf_ram.memory[4][3] ),
    .I1(\u_cpu.rf_ram.memory[5][3] ),
    .I2(\u_cpu.rf_ram.memory[6][3] ),
    .I3(\u_cpu.rf_ram.memory[7][3] ),
    .S0(_01959_),
    .S1(_02071_),
    .Z(_02072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06459_ (.A1(_01958_),
    .A2(_02072_),
    .ZN(_02073_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06460_ (.I(_01582_),
    .Z(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06461_ (.I0(\u_cpu.rf_ram.memory[0][3] ),
    .I1(\u_cpu.rf_ram.memory[1][3] ),
    .I2(\u_cpu.rf_ram.memory[2][3] ),
    .I3(\u_cpu.rf_ram.memory[3][3] ),
    .S0(_02074_),
    .S1(_01599_),
    .Z(_02075_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06462_ (.A1(_01597_),
    .A2(_02075_),
    .B(_01603_),
    .ZN(_02076_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06463_ (.A1(_02067_),
    .A2(_02070_),
    .B1(_02073_),
    .B2(_02076_),
    .C(_01607_),
    .ZN(_02077_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06464_ (.I(_01610_),
    .Z(_02078_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06465_ (.I0(\u_cpu.rf_ram.memory[20][3] ),
    .I1(\u_cpu.rf_ram.memory[21][3] ),
    .I2(\u_cpu.rf_ram.memory[22][3] ),
    .I3(\u_cpu.rf_ram.memory[23][3] ),
    .S0(_01849_),
    .S1(_01965_),
    .Z(_02079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06466_ (.A1(_02078_),
    .A2(_02079_),
    .ZN(_02080_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06467_ (.I(_01596_),
    .Z(_02081_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06468_ (.I0(\u_cpu.rf_ram.memory[16][3] ),
    .I1(\u_cpu.rf_ram.memory[17][3] ),
    .I2(\u_cpu.rf_ram.memory[18][3] ),
    .I3(\u_cpu.rf_ram.memory[19][3] ),
    .S0(_01852_),
    .S1(_01968_),
    .Z(_02082_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06469_ (.A1(_02081_),
    .A2(_02082_),
    .B(_01970_),
    .ZN(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06470_ (.I(_01573_),
    .Z(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06471_ (.I0(\u_cpu.rf_ram.memory[28][3] ),
    .I1(\u_cpu.rf_ram.memory[29][3] ),
    .I2(\u_cpu.rf_ram.memory[30][3] ),
    .I3(\u_cpu.rf_ram.memory[31][3] ),
    .S0(_02084_),
    .S1(_01634_),
    .Z(_02085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06472_ (.A1(_01630_),
    .A2(_02085_),
    .ZN(_02086_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06473_ (.I0(\u_cpu.rf_ram.memory[24][3] ),
    .I1(\u_cpu.rf_ram.memory[25][3] ),
    .I2(\u_cpu.rf_ram.memory[26][3] ),
    .I3(\u_cpu.rf_ram.memory[27][3] ),
    .S0(_01640_),
    .S1(_01642_),
    .Z(_02087_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06474_ (.A1(_01857_),
    .A2(_02087_),
    .B(_01859_),
    .ZN(_02088_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06475_ (.A1(_02080_),
    .A2(_02083_),
    .B1(_02086_),
    .B2(_02088_),
    .C(_01428_),
    .ZN(_02089_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06476_ (.I0(\u_cpu.rf_ram.memory[52][3] ),
    .I1(\u_cpu.rf_ram.memory[53][3] ),
    .I2(\u_cpu.rf_ram.memory[54][3] ),
    .I3(\u_cpu.rf_ram.memory[55][3] ),
    .S0(_01863_),
    .S1(_01653_),
    .Z(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06477_ (.A1(_01649_),
    .A2(_02090_),
    .ZN(_02091_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06478_ (.I(_01659_),
    .Z(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06479_ (.I0(\u_cpu.rf_ram.memory[48][3] ),
    .I1(\u_cpu.rf_ram.memory[49][3] ),
    .I2(\u_cpu.rf_ram.memory[50][3] ),
    .I3(\u_cpu.rf_ram.memory[51][3] ),
    .S0(_01657_),
    .S1(_02092_),
    .Z(_02093_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06480_ (.A1(_01656_),
    .A2(_02093_),
    .B(_01867_),
    .ZN(_02094_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06481_ (.I(_01638_),
    .Z(_02095_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06482_ (.I0(\u_cpu.rf_ram.memory[60][3] ),
    .I1(\u_cpu.rf_ram.memory[61][3] ),
    .I2(\u_cpu.rf_ram.memory[62][3] ),
    .I3(\u_cpu.rf_ram.memory[63][3] ),
    .S0(_02095_),
    .S1(_01668_),
    .Z(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06483_ (.A1(_01666_),
    .A2(_02096_),
    .ZN(_02097_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06484_ (.I(_01671_),
    .Z(_02098_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06485_ (.I(_01675_),
    .Z(_02099_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06486_ (.I0(\u_cpu.rf_ram.memory[56][3] ),
    .I1(\u_cpu.rf_ram.memory[57][3] ),
    .I2(\u_cpu.rf_ram.memory[58][3] ),
    .I3(\u_cpu.rf_ram.memory[59][3] ),
    .S0(_01871_),
    .S1(_02099_),
    .Z(_02100_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06487_ (.A1(_02098_),
    .A2(_02100_),
    .B(_01873_),
    .ZN(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06488_ (.A1(_02091_),
    .A2(_02094_),
    .B1(_02097_),
    .B2(_02101_),
    .C(_01681_),
    .ZN(_02102_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06489_ (.I(_01687_),
    .Z(_02103_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06490_ (.I0(\u_cpu.rf_ram.memory[40][3] ),
    .I1(\u_cpu.rf_ram.memory[41][3] ),
    .I2(\u_cpu.rf_ram.memory[42][3] ),
    .I3(\u_cpu.rf_ram.memory[43][3] ),
    .S0(_01686_),
    .S1(_02103_),
    .Z(_02104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06491_ (.A1(_01876_),
    .A2(_02104_),
    .ZN(_02105_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06492_ (.I0(\u_cpu.rf_ram.memory[44][3] ),
    .I1(\u_cpu.rf_ram.memory[45][3] ),
    .I2(\u_cpu.rf_ram.memory[46][3] ),
    .I3(\u_cpu.rf_ram.memory[47][3] ),
    .S0(_01692_),
    .S1(_01879_),
    .Z(_02106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06493_ (.I(_01417_),
    .Z(_02107_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06494_ (.A1(_01988_),
    .A2(_02106_),
    .B(_02107_),
    .ZN(_02108_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06495_ (.I(_01667_),
    .Z(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06496_ (.I0(\u_cpu.rf_ram.memory[36][3] ),
    .I1(\u_cpu.rf_ram.memory[37][3] ),
    .I2(\u_cpu.rf_ram.memory[38][3] ),
    .I3(\u_cpu.rf_ram.memory[39][3] ),
    .S0(_01698_),
    .S1(_02109_),
    .Z(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06497_ (.A1(_01882_),
    .A2(_02110_),
    .ZN(_02111_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06498_ (.I0(\u_cpu.rf_ram.memory[32][3] ),
    .I1(\u_cpu.rf_ram.memory[33][3] ),
    .I2(\u_cpu.rf_ram.memory[34][3] ),
    .I3(\u_cpu.rf_ram.memory[35][3] ),
    .S0(_01705_),
    .S1(_01994_),
    .Z(_02112_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06499_ (.A1(_01993_),
    .A2(_02112_),
    .B(_01996_),
    .ZN(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06500_ (.A1(_02105_),
    .A2(_02108_),
    .B1(_02111_),
    .B2(_02113_),
    .C(_01711_),
    .ZN(_02114_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06501_ (.A1(_01862_),
    .A2(_02102_),
    .A3(_02114_),
    .Z(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06502_ (.A1(_01566_),
    .A2(_02077_),
    .A3(_02089_),
    .B(_02115_),
    .ZN(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06503_ (.I(_01665_),
    .Z(_02117_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06504_ (.I0(\u_cpu.rf_ram.memory[108][3] ),
    .I1(\u_cpu.rf_ram.memory[109][3] ),
    .I2(\u_cpu.rf_ram.memory[110][3] ),
    .I3(\u_cpu.rf_ram.memory[111][3] ),
    .S0(_02001_),
    .S1(_01717_),
    .Z(_02118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06505_ (.A1(_02117_),
    .A2(_02118_),
    .ZN(_02119_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06506_ (.I0(\u_cpu.rf_ram.memory[104][3] ),
    .I1(\u_cpu.rf_ram.memory[105][3] ),
    .I2(\u_cpu.rf_ram.memory[106][3] ),
    .I3(\u_cpu.rf_ram.memory[107][3] ),
    .S0(_02005_),
    .S1(_01892_),
    .Z(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06507_ (.A1(_02004_),
    .A2(_02120_),
    .B(_01723_),
    .ZN(_02121_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06508_ (.I(_01638_),
    .Z(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06509_ (.I0(\u_cpu.rf_ram.memory[100][3] ),
    .I1(\u_cpu.rf_ram.memory[101][3] ),
    .I2(\u_cpu.rf_ram.memory[102][3] ),
    .I3(\u_cpu.rf_ram.memory[103][3] ),
    .S0(_02122_),
    .S1(_01895_),
    .Z(_02123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06510_ (.A1(_02008_),
    .A2(_02123_),
    .ZN(_02124_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06511_ (.I(_01673_),
    .Z(_02125_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06512_ (.I0(\u_cpu.rf_ram.memory[96][3] ),
    .I1(\u_cpu.rf_ram.memory[97][3] ),
    .I2(\u_cpu.rf_ram.memory[98][3] ),
    .I3(\u_cpu.rf_ram.memory[99][3] ),
    .S0(_02125_),
    .S1(_01641_),
    .Z(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06513_ (.A1(_01728_),
    .A2(_02126_),
    .B(_01731_),
    .ZN(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06514_ (.A1(_02119_),
    .A2(_02121_),
    .B1(_02124_),
    .B2(_02127_),
    .C(_01900_),
    .ZN(_02128_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06515_ (.I0(\u_cpu.rf_ram.memory[124][3] ),
    .I1(\u_cpu.rf_ram.memory[125][3] ),
    .I2(\u_cpu.rf_ram.memory[126][3] ),
    .I3(\u_cpu.rf_ram.memory[127][3] ),
    .S0(_02015_),
    .S1(_01737_),
    .Z(_02129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06516_ (.A1(_02014_),
    .A2(_02129_),
    .ZN(_02130_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06517_ (.I0(\u_cpu.rf_ram.memory[120][3] ),
    .I1(\u_cpu.rf_ram.memory[121][3] ),
    .I2(\u_cpu.rf_ram.memory[122][3] ),
    .I3(\u_cpu.rf_ram.memory[123][3] ),
    .S0(_01741_),
    .S1(_01905_),
    .Z(_02131_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06518_ (.A1(_01904_),
    .A2(_02131_),
    .B(_01744_),
    .ZN(_02132_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06519_ (.I(_01650_),
    .Z(_02133_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06520_ (.I0(\u_cpu.rf_ram.memory[112][3] ),
    .I1(\u_cpu.rf_ram.memory[113][3] ),
    .I2(\u_cpu.rf_ram.memory[114][3] ),
    .I3(\u_cpu.rf_ram.memory[115][3] ),
    .S0(_02133_),
    .S1(_01908_),
    .Z(_02134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06521_ (.A1(_01746_),
    .A2(_02134_),
    .ZN(_02135_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06522_ (.I(_01704_),
    .Z(_02136_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06523_ (.I0(\u_cpu.rf_ram.memory[116][3] ),
    .I1(\u_cpu.rf_ram.memory[117][3] ),
    .I2(\u_cpu.rf_ram.memory[118][3] ),
    .I3(\u_cpu.rf_ram.memory[119][3] ),
    .S0(_02136_),
    .S1(_01753_),
    .Z(_02137_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06524_ (.A1(_01751_),
    .A2(_02137_),
    .B(_01755_),
    .ZN(_02138_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06525_ (.I(_01426_),
    .Z(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06526_ (.A1(_02130_),
    .A2(_02132_),
    .B1(_02135_),
    .B2(_02138_),
    .C(_02139_),
    .ZN(_02140_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06527_ (.A1(_01423_),
    .A2(_02128_),
    .A3(_02140_),
    .ZN(_02141_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06528_ (.I(_01685_),
    .Z(_02142_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06529_ (.I0(\u_cpu.rf_ram.memory[92][3] ),
    .I1(\u_cpu.rf_ram.memory[93][3] ),
    .I2(\u_cpu.rf_ram.memory[94][3] ),
    .I3(\u_cpu.rf_ram.memory[95][3] ),
    .S0(_02142_),
    .S1(_01915_),
    .Z(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06530_ (.A1(_01761_),
    .A2(_02143_),
    .ZN(_02144_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06531_ (.I0(\u_cpu.rf_ram.memory[88][3] ),
    .I1(\u_cpu.rf_ram.memory[89][3] ),
    .I2(\u_cpu.rf_ram.memory[90][3] ),
    .I3(\u_cpu.rf_ram.memory[91][3] ),
    .S0(_02029_),
    .S1(_01768_),
    .Z(_02145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06532_ (.A1(_01766_),
    .A2(_02145_),
    .B(_02031_),
    .ZN(_02146_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06533_ (.I(_01702_),
    .Z(_02147_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06534_ (.I0(\u_cpu.rf_ram.memory[80][3] ),
    .I1(\u_cpu.rf_ram.memory[81][3] ),
    .I2(\u_cpu.rf_ram.memory[82][3] ),
    .I3(\u_cpu.rf_ram.memory[83][3] ),
    .S0(_01773_),
    .S1(_02033_),
    .Z(_02148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06535_ (.A1(_02147_),
    .A2(_02148_),
    .ZN(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06536_ (.I(_01609_),
    .Z(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06537_ (.I(_01632_),
    .Z(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06538_ (.I0(\u_cpu.rf_ram.memory[84][3] ),
    .I1(\u_cpu.rf_ram.memory[85][3] ),
    .I2(\u_cpu.rf_ram.memory[86][3] ),
    .I3(\u_cpu.rf_ram.memory[87][3] ),
    .S0(_01922_),
    .S1(_02151_),
    .Z(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06539_ (.I(_01627_),
    .Z(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06540_ (.A1(_02150_),
    .A2(_02152_),
    .B(_02153_),
    .ZN(_02154_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06541_ (.A1(_02144_),
    .A2(_02146_),
    .B1(_02149_),
    .B2(_02154_),
    .C(_01925_),
    .ZN(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06542_ (.I0(\u_cpu.rf_ram.memory[64][3] ),
    .I1(\u_cpu.rf_ram.memory[65][3] ),
    .I2(\u_cpu.rf_ram.memory[66][3] ),
    .I3(\u_cpu.rf_ram.memory[67][3] ),
    .S0(_01787_),
    .S1(_02040_),
    .Z(_02156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06543_ (.A1(_02039_),
    .A2(_02156_),
    .ZN(_02157_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06544_ (.I0(\u_cpu.rf_ram.memory[68][3] ),
    .I1(\u_cpu.rf_ram.memory[69][3] ),
    .I2(\u_cpu.rf_ram.memory[70][3] ),
    .I3(\u_cpu.rf_ram.memory[71][3] ),
    .S0(_01792_),
    .S1(_01930_),
    .Z(_02158_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06545_ (.A1(_01929_),
    .A2(_02158_),
    .B(_01932_),
    .ZN(_02159_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06546_ (.I0(\u_cpu.rf_ram.memory[72][3] ),
    .I1(\u_cpu.rf_ram.memory[73][3] ),
    .I2(\u_cpu.rf_ram.memory[74][3] ),
    .I3(\u_cpu.rf_ram.memory[75][3] ),
    .S0(_01934_),
    .S1(_01799_),
    .Z(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06547_ (.A1(_01797_),
    .A2(_02160_),
    .ZN(_02161_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06548_ (.I0(\u_cpu.rf_ram.memory[76][3] ),
    .I1(\u_cpu.rf_ram.memory[77][3] ),
    .I2(\u_cpu.rf_ram.memory[78][3] ),
    .I3(\u_cpu.rf_ram.memory[79][3] ),
    .S0(_02047_),
    .S1(_01803_),
    .Z(_02162_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06549_ (.A1(_01802_),
    .A2(_02162_),
    .B(_01805_),
    .ZN(_02163_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06550_ (.A1(_02157_),
    .A2(_02159_),
    .B1(_02161_),
    .B2(_02163_),
    .C(_02050_),
    .ZN(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06551_ (.A1(_02026_),
    .A2(_02155_),
    .A3(_02164_),
    .ZN(_02165_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06552_ (.A1(_02141_),
    .A2(_02165_),
    .B(_01810_),
    .ZN(_02166_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06553_ (.I0(\u_cpu.rf_ram.memory[136][3] ),
    .I1(\u_cpu.rf_ram.memory[137][3] ),
    .I2(\u_cpu.rf_ram.memory[138][3] ),
    .I3(\u_cpu.rf_ram.memory[139][3] ),
    .S0(_01814_),
    .S1(_01942_),
    .Z(_02167_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06554_ (.A1(_01400_),
    .A2(_02167_),
    .ZN(_02168_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06555_ (.I(_01813_),
    .Z(_02169_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06556_ (.I0(\u_cpu.rf_ram.memory[140][3] ),
    .I1(\u_cpu.rf_ram.memory[141][3] ),
    .I2(\u_cpu.rf_ram.memory[142][3] ),
    .I3(\u_cpu.rf_ram.memory[143][3] ),
    .S0(_02169_),
    .S1(_01821_),
    .Z(_02170_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06557_ (.A1(_01819_),
    .A2(_02170_),
    .B(_01823_),
    .ZN(_02171_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06558_ (.I0(\u_cpu.rf_ram.memory[128][3] ),
    .I1(\u_cpu.rf_ram.memory[129][3] ),
    .I2(\u_cpu.rf_ram.memory[130][3] ),
    .I3(\u_cpu.rf_ram.memory[131][3] ),
    .S0(_01826_),
    .S1(_01827_),
    .Z(_02172_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06559_ (.A1(_01947_),
    .A2(_02172_),
    .ZN(_02173_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06560_ (.I(_01788_),
    .Z(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06561_ (.I0(\u_cpu.rf_ram.memory[132][3] ),
    .I1(\u_cpu.rf_ram.memory[133][3] ),
    .I2(\u_cpu.rf_ram.memory[134][3] ),
    .I3(\u_cpu.rf_ram.memory[135][3] ),
    .S0(_02061_),
    .S1(_02174_),
    .Z(_02175_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06562_ (.A1(_02060_),
    .A2(_02175_),
    .B(_01419_),
    .ZN(_02176_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _06563_ (.A1(_02168_),
    .A2(_02171_),
    .B1(_02173_),
    .B2(_02176_),
    .C(_01835_),
    .ZN(_02177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06564_ (.A1(_02166_),
    .A2(_02177_),
    .ZN(_02178_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06565_ (.A1(_01564_),
    .A2(_02116_),
    .B(_02178_),
    .ZN(_00003_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06566_ (.I0(\u_cpu.rf_ram.memory[8][4] ),
    .I1(\u_cpu.rf_ram.memory[9][4] ),
    .I2(\u_cpu.rf_ram.memory[10][4] ),
    .I3(\u_cpu.rf_ram.memory[11][4] ),
    .S0(_01574_),
    .S1(_01838_),
    .Z(_02179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06567_ (.A1(_01637_),
    .A2(_02179_),
    .ZN(_02180_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06568_ (.I0(\u_cpu.rf_ram.memory[12][4] ),
    .I1(\u_cpu.rf_ram.memory[13][4] ),
    .I2(\u_cpu.rf_ram.memory[14][4] ),
    .I3(\u_cpu.rf_ram.memory[15][4] ),
    .S0(_01583_),
    .S1(_01841_),
    .Z(_02181_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06569_ (.A1(_01399_),
    .A2(_02181_),
    .B(_02069_),
    .ZN(_02182_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06570_ (.I0(\u_cpu.rf_ram.memory[4][4] ),
    .I1(\u_cpu.rf_ram.memory[5][4] ),
    .I2(\u_cpu.rf_ram.memory[6][4] ),
    .I3(\u_cpu.rf_ram.memory[7][4] ),
    .S0(_01959_),
    .S1(_02071_),
    .Z(_02183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06571_ (.A1(_01958_),
    .A2(_02183_),
    .ZN(_02184_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06572_ (.I0(\u_cpu.rf_ram.memory[0][4] ),
    .I1(\u_cpu.rf_ram.memory[1][4] ),
    .I2(\u_cpu.rf_ram.memory[2][4] ),
    .I3(\u_cpu.rf_ram.memory[3][4] ),
    .S0(_02074_),
    .S1(_01585_),
    .Z(_02185_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06573_ (.A1(_01597_),
    .A2(_02185_),
    .B(_01795_),
    .ZN(_02186_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06574_ (.A1(_02180_),
    .A2(_02182_),
    .B1(_02184_),
    .B2(_02186_),
    .C(_01607_),
    .ZN(_02187_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06575_ (.I0(\u_cpu.rf_ram.memory[20][4] ),
    .I1(\u_cpu.rf_ram.memory[21][4] ),
    .I2(\u_cpu.rf_ram.memory[22][4] ),
    .I3(\u_cpu.rf_ram.memory[23][4] ),
    .S0(_01849_),
    .S1(_01965_),
    .Z(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06576_ (.A1(_02078_),
    .A2(_02188_),
    .ZN(_02189_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06577_ (.I0(\u_cpu.rf_ram.memory[16][4] ),
    .I1(\u_cpu.rf_ram.memory[17][4] ),
    .I2(\u_cpu.rf_ram.memory[18][4] ),
    .I3(\u_cpu.rf_ram.memory[19][4] ),
    .S0(_01852_),
    .S1(_01968_),
    .Z(_02190_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06578_ (.A1(_02081_),
    .A2(_02190_),
    .B(_01970_),
    .ZN(_02191_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06579_ (.I0(\u_cpu.rf_ram.memory[28][4] ),
    .I1(\u_cpu.rf_ram.memory[29][4] ),
    .I2(\u_cpu.rf_ram.memory[30][4] ),
    .I3(\u_cpu.rf_ram.memory[31][4] ),
    .S0(_02084_),
    .S1(_01577_),
    .Z(_02192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06580_ (.A1(_01630_),
    .A2(_02192_),
    .ZN(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06581_ (.I0(\u_cpu.rf_ram.memory[24][4] ),
    .I1(\u_cpu.rf_ram.memory[25][4] ),
    .I2(\u_cpu.rf_ram.memory[26][4] ),
    .I3(\u_cpu.rf_ram.memory[27][4] ),
    .S0(_01622_),
    .S1(_01642_),
    .Z(_02194_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06582_ (.A1(_01857_),
    .A2(_02194_),
    .B(_01859_),
    .ZN(_02195_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06583_ (.A1(_02189_),
    .A2(_02191_),
    .B1(_02193_),
    .B2(_02195_),
    .C(_01784_),
    .ZN(_02196_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06584_ (.I0(\u_cpu.rf_ram.memory[52][4] ),
    .I1(\u_cpu.rf_ram.memory[53][4] ),
    .I2(\u_cpu.rf_ram.memory[54][4] ),
    .I3(\u_cpu.rf_ram.memory[55][4] ),
    .S0(_01863_),
    .S1(_01748_),
    .Z(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06585_ (.A1(_01697_),
    .A2(_02197_),
    .ZN(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06586_ (.I0(\u_cpu.rf_ram.memory[48][4] ),
    .I1(\u_cpu.rf_ram.memory[49][4] ),
    .I2(\u_cpu.rf_ram.memory[50][4] ),
    .I3(\u_cpu.rf_ram.memory[51][4] ),
    .S0(_01812_),
    .S1(_02092_),
    .Z(_02199_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06587_ (.A1(_01569_),
    .A2(_02199_),
    .B(_01867_),
    .ZN(_02200_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06588_ (.I0(\u_cpu.rf_ram.memory[60][4] ),
    .I1(\u_cpu.rf_ram.memory[61][4] ),
    .I2(\u_cpu.rf_ram.memory[62][4] ),
    .I3(\u_cpu.rf_ram.memory[63][4] ),
    .S0(_02095_),
    .S1(_01668_),
    .Z(_02201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06589_ (.A1(_01666_),
    .A2(_02201_),
    .ZN(_02202_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06590_ (.I0(\u_cpu.rf_ram.memory[56][4] ),
    .I1(\u_cpu.rf_ram.memory[57][4] ),
    .I2(\u_cpu.rf_ram.memory[58][4] ),
    .I3(\u_cpu.rf_ram.memory[59][4] ),
    .S0(_01871_),
    .S1(_02099_),
    .Z(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06591_ (.A1(_02098_),
    .A2(_02203_),
    .B(_01873_),
    .ZN(_02204_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06592_ (.A1(_02198_),
    .A2(_02200_),
    .B1(_02202_),
    .B2(_02204_),
    .C(_01681_),
    .ZN(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06593_ (.I0(\u_cpu.rf_ram.memory[40][4] ),
    .I1(\u_cpu.rf_ram.memory[41][4] ),
    .I2(\u_cpu.rf_ram.memory[42][4] ),
    .I3(\u_cpu.rf_ram.memory[43][4] ),
    .S0(_01686_),
    .S1(_02103_),
    .Z(_02206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06594_ (.A1(_01876_),
    .A2(_02206_),
    .ZN(_02207_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06595_ (.I0(\u_cpu.rf_ram.memory[44][4] ),
    .I1(\u_cpu.rf_ram.memory[45][4] ),
    .I2(\u_cpu.rf_ram.memory[46][4] ),
    .I3(\u_cpu.rf_ram.memory[47][4] ),
    .S0(_01692_),
    .S1(_01879_),
    .Z(_02208_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06596_ (.A1(_01988_),
    .A2(_02208_),
    .B(_02107_),
    .ZN(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06597_ (.I0(\u_cpu.rf_ram.memory[36][4] ),
    .I1(\u_cpu.rf_ram.memory[37][4] ),
    .I2(\u_cpu.rf_ram.memory[38][4] ),
    .I3(\u_cpu.rf_ram.memory[39][4] ),
    .S0(_01698_),
    .S1(_02109_),
    .Z(_02210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06598_ (.A1(_01882_),
    .A2(_02210_),
    .ZN(_02211_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06599_ (.I0(\u_cpu.rf_ram.memory[32][4] ),
    .I1(\u_cpu.rf_ram.memory[33][4] ),
    .I2(\u_cpu.rf_ram.memory[34][4] ),
    .I3(\u_cpu.rf_ram.memory[35][4] ),
    .S0(_01705_),
    .S1(_01994_),
    .Z(_02212_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06600_ (.A1(_01993_),
    .A2(_02212_),
    .B(_01996_),
    .ZN(_02213_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06601_ (.A1(_02207_),
    .A2(_02209_),
    .B1(_02211_),
    .B2(_02213_),
    .C(_01733_),
    .ZN(_02214_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06602_ (.A1(_01862_),
    .A2(_02205_),
    .A3(_02214_),
    .Z(_02215_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06603_ (.A1(_01566_),
    .A2(_02187_),
    .A3(_02196_),
    .B(_02215_),
    .ZN(_02216_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06604_ (.I0(\u_cpu.rf_ram.memory[108][4] ),
    .I1(\u_cpu.rf_ram.memory[109][4] ),
    .I2(\u_cpu.rf_ram.memory[110][4] ),
    .I3(\u_cpu.rf_ram.memory[111][4] ),
    .S0(_02001_),
    .S1(_01717_),
    .Z(_02217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06605_ (.A1(_02117_),
    .A2(_02217_),
    .ZN(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06606_ (.I0(\u_cpu.rf_ram.memory[104][4] ),
    .I1(\u_cpu.rf_ram.memory[105][4] ),
    .I2(\u_cpu.rf_ram.memory[106][4] ),
    .I3(\u_cpu.rf_ram.memory[107][4] ),
    .S0(_02005_),
    .S1(_01892_),
    .Z(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06607_ (.A1(_02004_),
    .A2(_02219_),
    .B(_01723_),
    .ZN(_02220_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06608_ (.I0(\u_cpu.rf_ram.memory[100][4] ),
    .I1(\u_cpu.rf_ram.memory[101][4] ),
    .I2(\u_cpu.rf_ram.memory[102][4] ),
    .I3(\u_cpu.rf_ram.memory[103][4] ),
    .S0(_02122_),
    .S1(_01895_),
    .Z(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06609_ (.A1(_02008_),
    .A2(_02221_),
    .ZN(_02222_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06610_ (.I0(\u_cpu.rf_ram.memory[96][4] ),
    .I1(\u_cpu.rf_ram.memory[97][4] ),
    .I2(\u_cpu.rf_ram.memory[98][4] ),
    .I3(\u_cpu.rf_ram.memory[99][4] ),
    .S0(_02125_),
    .S1(_01693_),
    .Z(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06611_ (.A1(_01728_),
    .A2(_02223_),
    .B(_01663_),
    .ZN(_02224_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06612_ (.A1(_02218_),
    .A2(_02220_),
    .B1(_02222_),
    .B2(_02224_),
    .C(_01900_),
    .ZN(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06613_ (.I0(\u_cpu.rf_ram.memory[124][4] ),
    .I1(\u_cpu.rf_ram.memory[125][4] ),
    .I2(\u_cpu.rf_ram.memory[126][4] ),
    .I3(\u_cpu.rf_ram.memory[127][4] ),
    .S0(_02015_),
    .S1(_01737_),
    .Z(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06614_ (.A1(_02014_),
    .A2(_02226_),
    .ZN(_02227_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06615_ (.I0(\u_cpu.rf_ram.memory[120][4] ),
    .I1(\u_cpu.rf_ram.memory[121][4] ),
    .I2(\u_cpu.rf_ram.memory[122][4] ),
    .I3(\u_cpu.rf_ram.memory[123][4] ),
    .S0(_01674_),
    .S1(_01905_),
    .Z(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06616_ (.A1(_01904_),
    .A2(_02228_),
    .B(_01679_),
    .ZN(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06617_ (.I0(\u_cpu.rf_ram.memory[112][4] ),
    .I1(\u_cpu.rf_ram.memory[113][4] ),
    .I2(\u_cpu.rf_ram.memory[114][4] ),
    .I3(\u_cpu.rf_ram.memory[115][4] ),
    .S0(_02133_),
    .S1(_01908_),
    .Z(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06618_ (.A1(_01746_),
    .A2(_02230_),
    .ZN(_02231_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06619_ (.I0(\u_cpu.rf_ram.memory[116][4] ),
    .I1(\u_cpu.rf_ram.memory[117][4] ),
    .I2(\u_cpu.rf_ram.memory[118][4] ),
    .I3(\u_cpu.rf_ram.memory[119][4] ),
    .S0(_02136_),
    .S1(_01753_),
    .Z(_02232_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06620_ (.A1(_01751_),
    .A2(_02232_),
    .B(_01755_),
    .ZN(_02233_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06621_ (.A1(_02227_),
    .A2(_02229_),
    .B1(_02231_),
    .B2(_02233_),
    .C(_02139_),
    .ZN(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06622_ (.A1(_01647_),
    .A2(_02225_),
    .A3(_02234_),
    .ZN(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06623_ (.I0(\u_cpu.rf_ram.memory[92][4] ),
    .I1(\u_cpu.rf_ram.memory[93][4] ),
    .I2(\u_cpu.rf_ram.memory[94][4] ),
    .I3(\u_cpu.rf_ram.memory[95][4] ),
    .S0(_02142_),
    .S1(_01915_),
    .Z(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06624_ (.A1(_01761_),
    .A2(_02236_),
    .ZN(_02237_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06625_ (.I0(\u_cpu.rf_ram.memory[88][4] ),
    .I1(\u_cpu.rf_ram.memory[89][4] ),
    .I2(\u_cpu.rf_ram.memory[90][4] ),
    .I3(\u_cpu.rf_ram.memory[91][4] ),
    .S0(_02029_),
    .S1(_01742_),
    .Z(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06626_ (.A1(_01740_),
    .A2(_02238_),
    .B(_02031_),
    .ZN(_02239_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06627_ (.I0(\u_cpu.rf_ram.memory[80][4] ),
    .I1(\u_cpu.rf_ram.memory[81][4] ),
    .I2(\u_cpu.rf_ram.memory[82][4] ),
    .I3(\u_cpu.rf_ram.memory[83][4] ),
    .S0(_01651_),
    .S1(_02033_),
    .Z(_02240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06628_ (.A1(_02147_),
    .A2(_02240_),
    .ZN(_02241_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06629_ (.I0(\u_cpu.rf_ram.memory[84][4] ),
    .I1(\u_cpu.rf_ram.memory[85][4] ),
    .I2(\u_cpu.rf_ram.memory[86][4] ),
    .I3(\u_cpu.rf_ram.memory[87][4] ),
    .S0(_01922_),
    .S1(_02151_),
    .Z(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06630_ (.A1(_02150_),
    .A2(_02242_),
    .B(_02153_),
    .ZN(_02243_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06631_ (.A1(_02237_),
    .A2(_02239_),
    .B1(_02241_),
    .B2(_02243_),
    .C(_01925_),
    .ZN(_02244_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06632_ (.I0(\u_cpu.rf_ram.memory[64][4] ),
    .I1(\u_cpu.rf_ram.memory[65][4] ),
    .I2(\u_cpu.rf_ram.memory[66][4] ),
    .I3(\u_cpu.rf_ram.memory[67][4] ),
    .S0(_01798_),
    .S1(_02040_),
    .Z(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06633_ (.A1(_02039_),
    .A2(_02245_),
    .ZN(_02246_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06634_ (.I0(\u_cpu.rf_ram.memory[68][4] ),
    .I1(\u_cpu.rf_ram.memory[69][4] ),
    .I2(\u_cpu.rf_ram.memory[70][4] ),
    .I3(\u_cpu.rf_ram.memory[71][4] ),
    .S0(_01779_),
    .S1(_01930_),
    .Z(_02247_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06635_ (.A1(_01929_),
    .A2(_02247_),
    .B(_01932_),
    .ZN(_02248_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06636_ (.I0(\u_cpu.rf_ram.memory[72][4] ),
    .I1(\u_cpu.rf_ram.memory[73][4] ),
    .I2(\u_cpu.rf_ram.memory[74][4] ),
    .I3(\u_cpu.rf_ram.memory[75][4] ),
    .S0(_01934_),
    .S1(_01763_),
    .Z(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06637_ (.A1(_01684_),
    .A2(_02249_),
    .ZN(_02250_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06638_ (.I0(\u_cpu.rf_ram.memory[76][4] ),
    .I1(\u_cpu.rf_ram.memory[77][4] ),
    .I2(\u_cpu.rf_ram.memory[78][4] ),
    .I3(\u_cpu.rf_ram.memory[79][4] ),
    .S0(_02047_),
    .S1(_01793_),
    .Z(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06639_ (.A1(_01791_),
    .A2(_02251_),
    .B(_01805_),
    .ZN(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06640_ (.A1(_02246_),
    .A2(_02248_),
    .B1(_02250_),
    .B2(_02252_),
    .C(_02050_),
    .ZN(_02253_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06641_ (.A1(_02026_),
    .A2(_02244_),
    .A3(_02253_),
    .ZN(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06642_ (.A1(_02235_),
    .A2(_02254_),
    .B(_01810_),
    .ZN(_02255_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06643_ (.I0(\u_cpu.rf_ram.memory[136][4] ),
    .I1(\u_cpu.rf_ram.memory[137][4] ),
    .I2(\u_cpu.rf_ram.memory[138][4] ),
    .I3(\u_cpu.rf_ram.memory[139][4] ),
    .S0(_01814_),
    .S1(_01942_),
    .Z(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06644_ (.A1(_01825_),
    .A2(_02256_),
    .ZN(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06645_ (.I0(\u_cpu.rf_ram.memory[140][4] ),
    .I1(\u_cpu.rf_ram.memory[141][4] ),
    .I2(\u_cpu.rf_ram.memory[142][4] ),
    .I3(\u_cpu.rf_ram.memory[143][4] ),
    .S0(_02169_),
    .S1(_01816_),
    .Z(_02258_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06646_ (.A1(_01819_),
    .A2(_02258_),
    .B(_01823_),
    .ZN(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06647_ (.I0(\u_cpu.rf_ram.memory[128][4] ),
    .I1(\u_cpu.rf_ram.memory[129][4] ),
    .I2(\u_cpu.rf_ram.memory[130][4] ),
    .I3(\u_cpu.rf_ram.memory[131][4] ),
    .S0(_01614_),
    .S1(_01827_),
    .Z(_02260_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06648_ (.A1(_01947_),
    .A2(_02260_),
    .ZN(_02261_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06649_ (.I0(\u_cpu.rf_ram.memory[132][4] ),
    .I1(\u_cpu.rf_ram.memory[133][4] ),
    .I2(\u_cpu.rf_ram.memory[134][4] ),
    .I3(\u_cpu.rf_ram.memory[135][4] ),
    .S0(_02061_),
    .S1(_02174_),
    .Z(_02262_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06650_ (.A1(_02060_),
    .A2(_02262_),
    .B(_01644_),
    .ZN(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _06651_ (.A1(_02257_),
    .A2(_02259_),
    .B1(_02261_),
    .B2(_02263_),
    .C(_01835_),
    .ZN(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06652_ (.A1(_02255_),
    .A2(_02264_),
    .ZN(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06653_ (.A1(_01564_),
    .A2(_02216_),
    .B(_02265_),
    .ZN(_00004_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06654_ (.I0(\u_cpu.rf_ram.memory[8][5] ),
    .I1(\u_cpu.rf_ram.memory[9][5] ),
    .I2(\u_cpu.rf_ram.memory[10][5] ),
    .I3(\u_cpu.rf_ram.memory[11][5] ),
    .S0(_01591_),
    .S1(_01838_),
    .Z(_02266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06655_ (.A1(_01637_),
    .A2(_02266_),
    .ZN(_02267_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06656_ (.I0(\u_cpu.rf_ram.memory[12][5] ),
    .I1(\u_cpu.rf_ram.memory[13][5] ),
    .I2(\u_cpu.rf_ram.memory[14][5] ),
    .I3(\u_cpu.rf_ram.memory[15][5] ),
    .S0(_01813_),
    .S1(_01841_),
    .Z(_02268_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06657_ (.A1(_01399_),
    .A2(_02268_),
    .B(_02069_),
    .ZN(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06658_ (.I0(\u_cpu.rf_ram.memory[4][5] ),
    .I1(\u_cpu.rf_ram.memory[5][5] ),
    .I2(\u_cpu.rf_ram.memory[6][5] ),
    .I3(\u_cpu.rf_ram.memory[7][5] ),
    .S0(_01959_),
    .S1(_02071_),
    .Z(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06659_ (.A1(_01958_),
    .A2(_02270_),
    .ZN(_02271_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06660_ (.I0(\u_cpu.rf_ram.memory[0][5] ),
    .I1(\u_cpu.rf_ram.memory[1][5] ),
    .I2(\u_cpu.rf_ram.memory[2][5] ),
    .I3(\u_cpu.rf_ram.memory[3][5] ),
    .S0(_02074_),
    .S1(_01585_),
    .Z(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06661_ (.A1(_01786_),
    .A2(_02272_),
    .B(_01795_),
    .ZN(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06662_ (.A1(_02267_),
    .A2(_02269_),
    .B1(_02271_),
    .B2(_02273_),
    .C(_01807_),
    .ZN(_02274_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06663_ (.I0(\u_cpu.rf_ram.memory[20][5] ),
    .I1(\u_cpu.rf_ram.memory[21][5] ),
    .I2(\u_cpu.rf_ram.memory[22][5] ),
    .I3(\u_cpu.rf_ram.memory[23][5] ),
    .S0(_01849_),
    .S1(_01965_),
    .Z(_02275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06664_ (.A1(_02078_),
    .A2(_02275_),
    .ZN(_02276_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06665_ (.I0(\u_cpu.rf_ram.memory[16][5] ),
    .I1(\u_cpu.rf_ram.memory[17][5] ),
    .I2(\u_cpu.rf_ram.memory[18][5] ),
    .I3(\u_cpu.rf_ram.memory[19][5] ),
    .S0(_01852_),
    .S1(_01968_),
    .Z(_02277_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06666_ (.A1(_02081_),
    .A2(_02277_),
    .B(_01970_),
    .ZN(_02278_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06667_ (.I0(\u_cpu.rf_ram.memory[28][5] ),
    .I1(\u_cpu.rf_ram.memory[29][5] ),
    .I2(\u_cpu.rf_ram.memory[30][5] ),
    .I3(\u_cpu.rf_ram.memory[31][5] ),
    .S0(_02084_),
    .S1(_01577_),
    .Z(_02279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06668_ (.A1(_01590_),
    .A2(_02279_),
    .ZN(_02280_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06669_ (.I0(\u_cpu.rf_ram.memory[24][5] ),
    .I1(\u_cpu.rf_ram.memory[25][5] ),
    .I2(\u_cpu.rf_ram.memory[26][5] ),
    .I3(\u_cpu.rf_ram.memory[27][5] ),
    .S0(_01622_),
    .S1(_01625_),
    .Z(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06670_ (.A1(_01857_),
    .A2(_02281_),
    .B(_01859_),
    .ZN(_02282_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06671_ (.A1(_02276_),
    .A2(_02278_),
    .B1(_02280_),
    .B2(_02282_),
    .C(_01784_),
    .ZN(_02283_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06672_ (.I0(\u_cpu.rf_ram.memory[52][5] ),
    .I1(\u_cpu.rf_ram.memory[53][5] ),
    .I2(\u_cpu.rf_ram.memory[54][5] ),
    .I3(\u_cpu.rf_ram.memory[55][5] ),
    .S0(_01863_),
    .S1(_01748_),
    .Z(_02284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06673_ (.A1(_01697_),
    .A2(_02284_),
    .ZN(_02285_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06674_ (.I0(\u_cpu.rf_ram.memory[48][5] ),
    .I1(\u_cpu.rf_ram.memory[49][5] ),
    .I2(\u_cpu.rf_ram.memory[50][5] ),
    .I3(\u_cpu.rf_ram.memory[51][5] ),
    .S0(_01812_),
    .S1(_02092_),
    .Z(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06675_ (.A1(_01569_),
    .A2(_02286_),
    .B(_01867_),
    .ZN(_02287_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06676_ (.I0(\u_cpu.rf_ram.memory[60][5] ),
    .I1(\u_cpu.rf_ram.memory[61][5] ),
    .I2(\u_cpu.rf_ram.memory[62][5] ),
    .I3(\u_cpu.rf_ram.memory[63][5] ),
    .S0(_02095_),
    .S1(_01633_),
    .Z(_02288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06677_ (.A1(_01725_),
    .A2(_02288_),
    .ZN(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06678_ (.I0(\u_cpu.rf_ram.memory[56][5] ),
    .I1(\u_cpu.rf_ram.memory[57][5] ),
    .I2(\u_cpu.rf_ram.memory[58][5] ),
    .I3(\u_cpu.rf_ram.memory[59][5] ),
    .S0(_01871_),
    .S1(_02099_),
    .Z(_02290_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06679_ (.A1(_02098_),
    .A2(_02290_),
    .B(_01873_),
    .ZN(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06680_ (.A1(_02285_),
    .A2(_02287_),
    .B1(_02289_),
    .B2(_02291_),
    .C(_01427_),
    .ZN(_02292_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06681_ (.I0(\u_cpu.rf_ram.memory[40][5] ),
    .I1(\u_cpu.rf_ram.memory[41][5] ),
    .I2(\u_cpu.rf_ram.memory[42][5] ),
    .I3(\u_cpu.rf_ram.memory[43][5] ),
    .S0(_01736_),
    .S1(_02103_),
    .Z(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06682_ (.A1(_01876_),
    .A2(_02293_),
    .ZN(_02294_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06683_ (.I0(\u_cpu.rf_ram.memory[44][5] ),
    .I1(\u_cpu.rf_ram.memory[45][5] ),
    .I2(\u_cpu.rf_ram.memory[46][5] ),
    .I3(\u_cpu.rf_ram.memory[47][5] ),
    .S0(_01721_),
    .S1(_01879_),
    .Z(_02295_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06684_ (.A1(_01988_),
    .A2(_02295_),
    .B(_02107_),
    .ZN(_02296_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06685_ (.I0(\u_cpu.rf_ram.memory[36][5] ),
    .I1(\u_cpu.rf_ram.memory[37][5] ),
    .I2(\u_cpu.rf_ram.memory[38][5] ),
    .I3(\u_cpu.rf_ram.memory[39][5] ),
    .S0(_01716_),
    .S1(_02109_),
    .Z(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06686_ (.A1(_01882_),
    .A2(_02297_),
    .ZN(_02298_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06687_ (.I0(\u_cpu.rf_ram.memory[32][5] ),
    .I1(\u_cpu.rf_ram.memory[33][5] ),
    .I2(\u_cpu.rf_ram.memory[34][5] ),
    .I3(\u_cpu.rf_ram.memory[35][5] ),
    .S0(_01767_),
    .S1(_01994_),
    .Z(_02299_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06688_ (.A1(_01993_),
    .A2(_02299_),
    .B(_01996_),
    .ZN(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06689_ (.A1(_02294_),
    .A2(_02296_),
    .B1(_02298_),
    .B2(_02300_),
    .C(_01733_),
    .ZN(_02301_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06690_ (.A1(_01862_),
    .A2(_02292_),
    .A3(_02301_),
    .Z(_02302_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06691_ (.A1(_01760_),
    .A2(_02274_),
    .A3(_02283_),
    .B(_02302_),
    .ZN(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06692_ (.I0(\u_cpu.rf_ram.memory[108][5] ),
    .I1(\u_cpu.rf_ram.memory[109][5] ),
    .I2(\u_cpu.rf_ram.memory[110][5] ),
    .I3(\u_cpu.rf_ram.memory[111][5] ),
    .S0(_02001_),
    .S1(_01615_),
    .Z(_02304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06693_ (.A1(_02117_),
    .A2(_02304_),
    .ZN(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06694_ (.I0(\u_cpu.rf_ram.memory[104][5] ),
    .I1(\u_cpu.rf_ram.memory[105][5] ),
    .I2(\u_cpu.rf_ram.memory[106][5] ),
    .I3(\u_cpu.rf_ram.memory[107][5] ),
    .S0(_02005_),
    .S1(_01892_),
    .Z(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06695_ (.A1(_02004_),
    .A2(_02306_),
    .B(_01587_),
    .ZN(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06696_ (.I0(\u_cpu.rf_ram.memory[100][5] ),
    .I1(\u_cpu.rf_ram.memory[101][5] ),
    .I2(\u_cpu.rf_ram.memory[102][5] ),
    .I3(\u_cpu.rf_ram.memory[103][5] ),
    .S0(_02122_),
    .S1(_01895_),
    .Z(_02308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06697_ (.A1(_02008_),
    .A2(_02308_),
    .ZN(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06698_ (.I0(\u_cpu.rf_ram.memory[96][5] ),
    .I1(\u_cpu.rf_ram.memory[97][5] ),
    .I2(\u_cpu.rf_ram.memory[98][5] ),
    .I3(\u_cpu.rf_ram.memory[99][5] ),
    .S0(_02125_),
    .S1(_01693_),
    .Z(_02310_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06699_ (.A1(_01720_),
    .A2(_02310_),
    .B(_01663_),
    .ZN(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06700_ (.A1(_02305_),
    .A2(_02307_),
    .B1(_02309_),
    .B2(_02311_),
    .C(_01900_),
    .ZN(_02312_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06701_ (.I0(\u_cpu.rf_ram.memory[124][5] ),
    .I1(\u_cpu.rf_ram.memory[125][5] ),
    .I2(\u_cpu.rf_ram.memory[126][5] ),
    .I3(\u_cpu.rf_ram.memory[127][5] ),
    .S0(_02015_),
    .S1(_01774_),
    .Z(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06702_ (.A1(_02014_),
    .A2(_02313_),
    .ZN(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06703_ (.I0(\u_cpu.rf_ram.memory[120][5] ),
    .I1(\u_cpu.rf_ram.memory[121][5] ),
    .I2(\u_cpu.rf_ram.memory[122][5] ),
    .I3(\u_cpu.rf_ram.memory[123][5] ),
    .S0(_01674_),
    .S1(_01905_),
    .Z(_02315_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06704_ (.A1(_01904_),
    .A2(_02315_),
    .B(_01679_),
    .ZN(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06705_ (.I0(\u_cpu.rf_ram.memory[112][5] ),
    .I1(\u_cpu.rf_ram.memory[113][5] ),
    .I2(\u_cpu.rf_ram.memory[114][5] ),
    .I3(\u_cpu.rf_ram.memory[115][5] ),
    .S0(_02133_),
    .S1(_01908_),
    .Z(_02317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06706_ (.A1(_01703_),
    .A2(_02317_),
    .ZN(_02318_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06707_ (.I0(\u_cpu.rf_ram.memory[116][5] ),
    .I1(\u_cpu.rf_ram.memory[117][5] ),
    .I2(\u_cpu.rf_ram.memory[118][5] ),
    .I3(\u_cpu.rf_ram.memory[119][5] ),
    .S0(_02136_),
    .S1(_01707_),
    .Z(_02319_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06708_ (.A1(_01691_),
    .A2(_02319_),
    .B(_01709_),
    .ZN(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06709_ (.A1(_02314_),
    .A2(_02316_),
    .B1(_02318_),
    .B2(_02320_),
    .C(_02139_),
    .ZN(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06710_ (.A1(_01647_),
    .A2(_02312_),
    .A3(_02321_),
    .ZN(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06711_ (.I0(\u_cpu.rf_ram.memory[92][5] ),
    .I1(\u_cpu.rf_ram.memory[93][5] ),
    .I2(\u_cpu.rf_ram.memory[94][5] ),
    .I3(\u_cpu.rf_ram.memory[95][5] ),
    .S0(_02142_),
    .S1(_01915_),
    .Z(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06712_ (.A1(_01735_),
    .A2(_02323_),
    .ZN(_02324_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06713_ (.I0(\u_cpu.rf_ram.memory[88][5] ),
    .I1(\u_cpu.rf_ram.memory[89][5] ),
    .I2(\u_cpu.rf_ram.memory[90][5] ),
    .I3(\u_cpu.rf_ram.memory[91][5] ),
    .S0(_02029_),
    .S1(_01742_),
    .Z(_02325_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06714_ (.A1(_01740_),
    .A2(_02325_),
    .B(_02031_),
    .ZN(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06715_ (.I0(\u_cpu.rf_ram.memory[80][5] ),
    .I1(\u_cpu.rf_ram.memory[81][5] ),
    .I2(\u_cpu.rf_ram.memory[82][5] ),
    .I3(\u_cpu.rf_ram.memory[83][5] ),
    .S0(_01651_),
    .S1(_02033_),
    .Z(_02327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06716_ (.A1(_02147_),
    .A2(_02327_),
    .ZN(_02328_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06717_ (.I0(\u_cpu.rf_ram.memory[84][5] ),
    .I1(\u_cpu.rf_ram.memory[85][5] ),
    .I2(\u_cpu.rf_ram.memory[86][5] ),
    .I3(\u_cpu.rf_ram.memory[87][5] ),
    .S0(_01922_),
    .S1(_02151_),
    .Z(_02329_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06718_ (.A1(_02150_),
    .A2(_02329_),
    .B(_02153_),
    .ZN(_02330_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06719_ (.A1(_02324_),
    .A2(_02326_),
    .B1(_02328_),
    .B2(_02330_),
    .C(_01925_),
    .ZN(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06720_ (.I0(\u_cpu.rf_ram.memory[64][5] ),
    .I1(\u_cpu.rf_ram.memory[65][5] ),
    .I2(\u_cpu.rf_ram.memory[66][5] ),
    .I3(\u_cpu.rf_ram.memory[67][5] ),
    .S0(_01798_),
    .S1(_02040_),
    .Z(_02332_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06721_ (.A1(_02039_),
    .A2(_02332_),
    .ZN(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06722_ (.I0(\u_cpu.rf_ram.memory[68][5] ),
    .I1(\u_cpu.rf_ram.memory[69][5] ),
    .I2(\u_cpu.rf_ram.memory[70][5] ),
    .I3(\u_cpu.rf_ram.memory[71][5] ),
    .S0(_01779_),
    .S1(_01930_),
    .Z(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06723_ (.A1(_01929_),
    .A2(_02334_),
    .B(_01932_),
    .ZN(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06724_ (.I0(\u_cpu.rf_ram.memory[72][5] ),
    .I1(\u_cpu.rf_ram.memory[73][5] ),
    .I2(\u_cpu.rf_ram.memory[74][5] ),
    .I3(\u_cpu.rf_ram.memory[75][5] ),
    .S0(_01934_),
    .S1(_01763_),
    .Z(_02336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06725_ (.A1(_01684_),
    .A2(_02336_),
    .ZN(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06726_ (.I0(\u_cpu.rf_ram.memory[76][5] ),
    .I1(\u_cpu.rf_ram.memory[77][5] ),
    .I2(\u_cpu.rf_ram.memory[78][5] ),
    .I3(\u_cpu.rf_ram.memory[79][5] ),
    .S0(_02047_),
    .S1(_01793_),
    .Z(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06727_ (.A1(_01791_),
    .A2(_02338_),
    .B(_01770_),
    .ZN(_02339_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06728_ (.A1(_02333_),
    .A2(_02335_),
    .B1(_02337_),
    .B2(_02339_),
    .C(_02050_),
    .ZN(_02340_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06729_ (.A1(_02026_),
    .A2(_02331_),
    .A3(_02340_),
    .ZN(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06730_ (.A1(_02322_),
    .A2(_02341_),
    .B(_01404_),
    .ZN(_02342_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06731_ (.I0(\u_cpu.rf_ram.memory[136][5] ),
    .I1(\u_cpu.rf_ram.memory[137][5] ),
    .I2(\u_cpu.rf_ram.memory[138][5] ),
    .I3(\u_cpu.rf_ram.memory[139][5] ),
    .S0(_01831_),
    .S1(_01942_),
    .Z(_02343_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06732_ (.A1(_01825_),
    .A2(_02343_),
    .ZN(_02344_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06733_ (.I0(\u_cpu.rf_ram.memory[140][5] ),
    .I1(\u_cpu.rf_ram.memory[141][5] ),
    .I2(\u_cpu.rf_ram.memory[142][5] ),
    .I3(\u_cpu.rf_ram.memory[143][5] ),
    .S0(_02169_),
    .S1(_01816_),
    .Z(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06734_ (.A1(_01830_),
    .A2(_02345_),
    .B(_01628_),
    .ZN(_02346_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06735_ (.I0(\u_cpu.rf_ram.memory[128][5] ),
    .I1(\u_cpu.rf_ram.memory[129][5] ),
    .I2(\u_cpu.rf_ram.memory[130][5] ),
    .I3(\u_cpu.rf_ram.memory[131][5] ),
    .S0(_01614_),
    .S1(_01616_),
    .Z(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06736_ (.A1(_01947_),
    .A2(_02347_),
    .ZN(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06737_ (.I0(\u_cpu.rf_ram.memory[132][5] ),
    .I1(\u_cpu.rf_ram.memory[133][5] ),
    .I2(\u_cpu.rf_ram.memory[134][5] ),
    .I3(\u_cpu.rf_ram.memory[135][5] ),
    .S0(_02061_),
    .S1(_02174_),
    .Z(_02349_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06738_ (.A1(_02060_),
    .A2(_02349_),
    .B(_01644_),
    .ZN(_02350_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _06739_ (.A1(_02344_),
    .A2(_02346_),
    .B1(_02348_),
    .B2(_02350_),
    .C(_01405_),
    .ZN(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06740_ (.A1(_02342_),
    .A2(_02351_),
    .ZN(_02352_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06741_ (.A1(_01406_),
    .A2(_02303_),
    .B(_02352_),
    .ZN(_00005_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06742_ (.I0(\u_cpu.rf_ram.memory[8][6] ),
    .I1(\u_cpu.rf_ram.memory[9][6] ),
    .I2(\u_cpu.rf_ram.memory[10][6] ),
    .I3(\u_cpu.rf_ram.memory[11][6] ),
    .S0(_01591_),
    .S1(_01592_),
    .Z(_02353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06743_ (.A1(_01637_),
    .A2(_02353_),
    .ZN(_02354_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06744_ (.I0(\u_cpu.rf_ram.memory[12][6] ),
    .I1(\u_cpu.rf_ram.memory[13][6] ),
    .I2(\u_cpu.rf_ram.memory[14][6] ),
    .I3(\u_cpu.rf_ram.memory[15][6] ),
    .S0(_01813_),
    .S1(_01815_),
    .Z(_02355_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06745_ (.A1(_01399_),
    .A2(_02355_),
    .B(_02069_),
    .ZN(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06746_ (.I0(\u_cpu.rf_ram.memory[4][6] ),
    .I1(\u_cpu.rf_ram.memory[5][6] ),
    .I2(\u_cpu.rf_ram.memory[6][6] ),
    .I3(\u_cpu.rf_ram.memory[7][6] ),
    .S0(_01959_),
    .S1(_02071_),
    .Z(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06747_ (.A1(_01958_),
    .A2(_02357_),
    .ZN(_02358_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06748_ (.I0(\u_cpu.rf_ram.memory[0][6] ),
    .I1(\u_cpu.rf_ram.memory[1][6] ),
    .I2(\u_cpu.rf_ram.memory[2][6] ),
    .I3(\u_cpu.rf_ram.memory[3][6] ),
    .S0(_02074_),
    .S1(_01585_),
    .Z(_02359_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06749_ (.A1(_01786_),
    .A2(_02359_),
    .B(_01795_),
    .ZN(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06750_ (.A1(_02354_),
    .A2(_02356_),
    .B1(_02358_),
    .B2(_02360_),
    .C(_01807_),
    .ZN(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06751_ (.I0(\u_cpu.rf_ram.memory[20][6] ),
    .I1(\u_cpu.rf_ram.memory[21][6] ),
    .I2(\u_cpu.rf_ram.memory[22][6] ),
    .I3(\u_cpu.rf_ram.memory[23][6] ),
    .S0(_01631_),
    .S1(_01965_),
    .Z(_02362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06752_ (.A1(_02078_),
    .A2(_02362_),
    .ZN(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06753_ (.I0(\u_cpu.rf_ram.memory[16][6] ),
    .I1(\u_cpu.rf_ram.memory[17][6] ),
    .I2(\u_cpu.rf_ram.memory[18][6] ),
    .I3(\u_cpu.rf_ram.memory[19][6] ),
    .S0(_01598_),
    .S1(_01968_),
    .Z(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06754_ (.A1(_02081_),
    .A2(_02364_),
    .B(_01970_),
    .ZN(_02365_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06755_ (.I0(\u_cpu.rf_ram.memory[28][6] ),
    .I1(\u_cpu.rf_ram.memory[29][6] ),
    .I2(\u_cpu.rf_ram.memory[30][6] ),
    .I3(\u_cpu.rf_ram.memory[31][6] ),
    .S0(_02084_),
    .S1(_01577_),
    .Z(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06756_ (.A1(_01590_),
    .A2(_02366_),
    .ZN(_02367_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06757_ (.I0(\u_cpu.rf_ram.memory[24][6] ),
    .I1(\u_cpu.rf_ram.memory[25][6] ),
    .I2(\u_cpu.rf_ram.memory[26][6] ),
    .I3(\u_cpu.rf_ram.memory[27][6] ),
    .S0(_01622_),
    .S1(_01625_),
    .Z(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06758_ (.A1(_01619_),
    .A2(_02368_),
    .B(_01588_),
    .ZN(_02369_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06759_ (.A1(_02363_),
    .A2(_02365_),
    .B1(_02367_),
    .B2(_02369_),
    .C(_01784_),
    .ZN(_02370_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06760_ (.I0(\u_cpu.rf_ram.memory[52][6] ),
    .I1(\u_cpu.rf_ram.memory[53][6] ),
    .I2(\u_cpu.rf_ram.memory[54][6] ),
    .I3(\u_cpu.rf_ram.memory[55][6] ),
    .S0(_01747_),
    .S1(_01748_),
    .Z(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06761_ (.A1(_01697_),
    .A2(_02371_),
    .ZN(_02372_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06762_ (.I0(\u_cpu.rf_ram.memory[48][6] ),
    .I1(\u_cpu.rf_ram.memory[49][6] ),
    .I2(\u_cpu.rf_ram.memory[50][6] ),
    .I3(\u_cpu.rf_ram.memory[51][6] ),
    .S0(_01812_),
    .S1(_02092_),
    .Z(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06763_ (.A1(_01569_),
    .A2(_02373_),
    .B(_01602_),
    .ZN(_02374_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06764_ (.I0(\u_cpu.rf_ram.memory[60][6] ),
    .I1(\u_cpu.rf_ram.memory[61][6] ),
    .I2(\u_cpu.rf_ram.memory[62][6] ),
    .I3(\u_cpu.rf_ram.memory[63][6] ),
    .S0(_02095_),
    .S1(_01633_),
    .Z(_02375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06765_ (.A1(_01725_),
    .A2(_02375_),
    .ZN(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06766_ (.I0(\u_cpu.rf_ram.memory[56][6] ),
    .I1(\u_cpu.rf_ram.memory[57][6] ),
    .I2(\u_cpu.rf_ram.memory[58][6] ),
    .I3(\u_cpu.rf_ram.memory[59][6] ),
    .S0(_01729_),
    .S1(_02099_),
    .Z(_02377_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06767_ (.A1(_02098_),
    .A2(_02377_),
    .B(_01695_),
    .ZN(_02378_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06768_ (.A1(_02372_),
    .A2(_02374_),
    .B1(_02376_),
    .B2(_02378_),
    .C(_01427_),
    .ZN(_02379_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06769_ (.I0(\u_cpu.rf_ram.memory[40][6] ),
    .I1(\u_cpu.rf_ram.memory[41][6] ),
    .I2(\u_cpu.rf_ram.memory[42][6] ),
    .I3(\u_cpu.rf_ram.memory[43][6] ),
    .S0(_01736_),
    .S1(_02103_),
    .Z(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06770_ (.A1(_01772_),
    .A2(_02380_),
    .ZN(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06771_ (.I0(\u_cpu.rf_ram.memory[44][6] ),
    .I1(\u_cpu.rf_ram.memory[45][6] ),
    .I2(\u_cpu.rf_ram.memory[46][6] ),
    .I3(\u_cpu.rf_ram.memory[47][6] ),
    .S0(_01721_),
    .S1(_01624_),
    .Z(_02382_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06772_ (.A1(_01988_),
    .A2(_02382_),
    .B(_02107_),
    .ZN(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06773_ (.I0(\u_cpu.rf_ram.memory[36][6] ),
    .I1(\u_cpu.rf_ram.memory[37][6] ),
    .I2(\u_cpu.rf_ram.memory[38][6] ),
    .I3(\u_cpu.rf_ram.memory[39][6] ),
    .S0(_01716_),
    .S1(_02109_),
    .Z(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06774_ (.A1(_01715_),
    .A2(_02384_),
    .ZN(_02385_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06775_ (.I0(\u_cpu.rf_ram.memory[32][6] ),
    .I1(\u_cpu.rf_ram.memory[33][6] ),
    .I2(\u_cpu.rf_ram.memory[34][6] ),
    .I3(\u_cpu.rf_ram.memory[35][6] ),
    .S0(_01767_),
    .S1(_01994_),
    .Z(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06776_ (.A1(_01993_),
    .A2(_02386_),
    .B(_01996_),
    .ZN(_02387_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06777_ (.A1(_02381_),
    .A2(_02383_),
    .B1(_02385_),
    .B2(_02387_),
    .C(_01733_),
    .ZN(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06778_ (.A1(_01422_),
    .A2(_02379_),
    .A3(_02388_),
    .Z(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06779_ (.A1(_01760_),
    .A2(_02361_),
    .A3(_02370_),
    .B(_02389_),
    .ZN(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06780_ (.I0(\u_cpu.rf_ram.memory[108][6] ),
    .I1(\u_cpu.rf_ram.memory[109][6] ),
    .I2(\u_cpu.rf_ram.memory[110][6] ),
    .I3(\u_cpu.rf_ram.memory[111][6] ),
    .S0(_02001_),
    .S1(_01615_),
    .Z(_02391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06781_ (.A1(_02117_),
    .A2(_02391_),
    .ZN(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06782_ (.I0(\u_cpu.rf_ram.memory[104][6] ),
    .I1(\u_cpu.rf_ram.memory[105][6] ),
    .I2(\u_cpu.rf_ram.memory[106][6] ),
    .I3(\u_cpu.rf_ram.memory[107][6] ),
    .S0(_02005_),
    .S1(_01660_),
    .Z(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06783_ (.A1(_02004_),
    .A2(_02393_),
    .B(_01587_),
    .ZN(_02394_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06784_ (.I0(\u_cpu.rf_ram.memory[100][6] ),
    .I1(\u_cpu.rf_ram.memory[101][6] ),
    .I2(\u_cpu.rf_ram.memory[102][6] ),
    .I3(\u_cpu.rf_ram.memory[103][6] ),
    .S0(_02122_),
    .S1(_01576_),
    .Z(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06785_ (.A1(_02008_),
    .A2(_02395_),
    .ZN(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06786_ (.I0(\u_cpu.rf_ram.memory[96][6] ),
    .I1(\u_cpu.rf_ram.memory[97][6] ),
    .I2(\u_cpu.rf_ram.memory[98][6] ),
    .I3(\u_cpu.rf_ram.memory[99][6] ),
    .S0(_02125_),
    .S1(_01693_),
    .Z(_02397_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06787_ (.A1(_01720_),
    .A2(_02397_),
    .B(_01663_),
    .ZN(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06788_ (.A1(_02392_),
    .A2(_02394_),
    .B1(_02396_),
    .B2(_02398_),
    .C(_01606_),
    .ZN(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06789_ (.I0(\u_cpu.rf_ram.memory[124][6] ),
    .I1(\u_cpu.rf_ram.memory[125][6] ),
    .I2(\u_cpu.rf_ram.memory[126][6] ),
    .I3(\u_cpu.rf_ram.memory[127][6] ),
    .S0(_02015_),
    .S1(_01774_),
    .Z(_02400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06790_ (.A1(_02014_),
    .A2(_02400_),
    .ZN(_02401_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06791_ (.I0(\u_cpu.rf_ram.memory[120][6] ),
    .I1(\u_cpu.rf_ram.memory[121][6] ),
    .I2(\u_cpu.rf_ram.memory[122][6] ),
    .I3(\u_cpu.rf_ram.memory[123][6] ),
    .S0(_01674_),
    .S1(_01676_),
    .Z(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06792_ (.A1(_01672_),
    .A2(_02402_),
    .B(_01679_),
    .ZN(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06793_ (.I0(\u_cpu.rf_ram.memory[112][6] ),
    .I1(\u_cpu.rf_ram.memory[113][6] ),
    .I2(\u_cpu.rf_ram.memory[114][6] ),
    .I3(\u_cpu.rf_ram.memory[115][6] ),
    .S0(_02133_),
    .S1(_01699_),
    .Z(_02404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06794_ (.A1(_01703_),
    .A2(_02404_),
    .ZN(_02405_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06795_ (.I0(\u_cpu.rf_ram.memory[116][6] ),
    .I1(\u_cpu.rf_ram.memory[117][6] ),
    .I2(\u_cpu.rf_ram.memory[118][6] ),
    .I3(\u_cpu.rf_ram.memory[119][6] ),
    .S0(_02136_),
    .S1(_01707_),
    .Z(_02406_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06796_ (.A1(_01691_),
    .A2(_02406_),
    .B(_01709_),
    .ZN(_02407_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06797_ (.A1(_02401_),
    .A2(_02403_),
    .B1(_02405_),
    .B2(_02407_),
    .C(_02139_),
    .ZN(_02408_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06798_ (.A1(_01647_),
    .A2(_02399_),
    .A3(_02408_),
    .ZN(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06799_ (.I0(\u_cpu.rf_ram.memory[92][6] ),
    .I1(\u_cpu.rf_ram.memory[93][6] ),
    .I2(\u_cpu.rf_ram.memory[94][6] ),
    .I3(\u_cpu.rf_ram.memory[95][6] ),
    .S0(_02142_),
    .S1(_01688_),
    .Z(_02410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06800_ (.A1(_01735_),
    .A2(_02410_),
    .ZN(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06801_ (.I0(\u_cpu.rf_ram.memory[88][6] ),
    .I1(\u_cpu.rf_ram.memory[89][6] ),
    .I2(\u_cpu.rf_ram.memory[90][6] ),
    .I3(\u_cpu.rf_ram.memory[91][6] ),
    .S0(_02029_),
    .S1(_01742_),
    .Z(_02412_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06802_ (.A1(_01740_),
    .A2(_02412_),
    .B(_02031_),
    .ZN(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06803_ (.I0(\u_cpu.rf_ram.memory[80][6] ),
    .I1(\u_cpu.rf_ram.memory[81][6] ),
    .I2(\u_cpu.rf_ram.memory[82][6] ),
    .I3(\u_cpu.rf_ram.memory[83][6] ),
    .S0(_01651_),
    .S1(_02033_),
    .Z(_02414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06804_ (.A1(_02147_),
    .A2(_02414_),
    .ZN(_02415_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06805_ (.I0(\u_cpu.rf_ram.memory[84][6] ),
    .I1(\u_cpu.rf_ram.memory[85][6] ),
    .I2(\u_cpu.rf_ram.memory[86][6] ),
    .I3(\u_cpu.rf_ram.memory[87][6] ),
    .S0(_01752_),
    .S1(_02151_),
    .Z(_02416_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06806_ (.A1(_02150_),
    .A2(_02416_),
    .B(_02153_),
    .ZN(_02417_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06807_ (.A1(_02411_),
    .A2(_02413_),
    .B1(_02415_),
    .B2(_02417_),
    .C(_01757_),
    .ZN(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06808_ (.I0(\u_cpu.rf_ram.memory[64][6] ),
    .I1(\u_cpu.rf_ram.memory[65][6] ),
    .I2(\u_cpu.rf_ram.memory[66][6] ),
    .I3(\u_cpu.rf_ram.memory[67][6] ),
    .S0(_01798_),
    .S1(_02040_),
    .Z(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06809_ (.A1(_02039_),
    .A2(_02419_),
    .ZN(_02420_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06810_ (.I0(\u_cpu.rf_ram.memory[68][6] ),
    .I1(\u_cpu.rf_ram.memory[69][6] ),
    .I2(\u_cpu.rf_ram.memory[70][6] ),
    .I3(\u_cpu.rf_ram.memory[71][6] ),
    .S0(_01779_),
    .S1(_01780_),
    .Z(_02421_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06811_ (.A1(_01778_),
    .A2(_02421_),
    .B(_01782_),
    .ZN(_02422_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06812_ (.I0(\u_cpu.rf_ram.memory[72][6] ),
    .I1(\u_cpu.rf_ram.memory[73][6] ),
    .I2(\u_cpu.rf_ram.memory[74][6] ),
    .I3(\u_cpu.rf_ram.memory[75][6] ),
    .S0(_01762_),
    .S1(_01763_),
    .Z(_02423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06813_ (.A1(_01684_),
    .A2(_02423_),
    .ZN(_02424_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06814_ (.I0(\u_cpu.rf_ram.memory[76][6] ),
    .I1(\u_cpu.rf_ram.memory[77][6] ),
    .I2(\u_cpu.rf_ram.memory[78][6] ),
    .I3(\u_cpu.rf_ram.memory[79][6] ),
    .S0(_02047_),
    .S1(_01793_),
    .Z(_02425_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06815_ (.A1(_01791_),
    .A2(_02425_),
    .B(_01770_),
    .ZN(_02426_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06816_ (.A1(_02420_),
    .A2(_02422_),
    .B1(_02424_),
    .B2(_02426_),
    .C(_02050_),
    .ZN(_02427_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06817_ (.A1(_02026_),
    .A2(_02418_),
    .A3(_02427_),
    .ZN(_02428_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06818_ (.A1(_02409_),
    .A2(_02428_),
    .B(_01404_),
    .ZN(_02429_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06819_ (.I0(\u_cpu.rf_ram.memory[136][6] ),
    .I1(\u_cpu.rf_ram.memory[137][6] ),
    .I2(\u_cpu.rf_ram.memory[138][6] ),
    .I3(\u_cpu.rf_ram.memory[139][6] ),
    .S0(_01831_),
    .S1(_01832_),
    .Z(_02430_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06820_ (.A1(_01825_),
    .A2(_02430_),
    .ZN(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06821_ (.I0(\u_cpu.rf_ram.memory[140][6] ),
    .I1(\u_cpu.rf_ram.memory[141][6] ),
    .I2(\u_cpu.rf_ram.memory[142][6] ),
    .I3(\u_cpu.rf_ram.memory[143][6] ),
    .S0(_02169_),
    .S1(_01816_),
    .Z(_02432_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06822_ (.A1(_01830_),
    .A2(_02432_),
    .B(_01628_),
    .ZN(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06823_ (.I0(\u_cpu.rf_ram.memory[128][6] ),
    .I1(\u_cpu.rf_ram.memory[129][6] ),
    .I2(\u_cpu.rf_ram.memory[130][6] ),
    .I3(\u_cpu.rf_ram.memory[131][6] ),
    .S0(_01614_),
    .S1(_01616_),
    .Z(_02434_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06824_ (.A1(_01611_),
    .A2(_02434_),
    .ZN(_02435_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06825_ (.I0(\u_cpu.rf_ram.memory[132][6] ),
    .I1(\u_cpu.rf_ram.memory[133][6] ),
    .I2(\u_cpu.rf_ram.memory[134][6] ),
    .I3(\u_cpu.rf_ram.memory[135][6] ),
    .S0(_02061_),
    .S1(_02174_),
    .Z(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06826_ (.A1(_02060_),
    .A2(_02436_),
    .B(_01644_),
    .ZN(_02437_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _06827_ (.A1(_02431_),
    .A2(_02433_),
    .B1(_02435_),
    .B2(_02437_),
    .C(_01405_),
    .ZN(_02438_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06828_ (.A1(_02429_),
    .A2(_02438_),
    .ZN(_02439_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06829_ (.A1(_01406_),
    .A2(_02390_),
    .B(_02439_),
    .ZN(_00006_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06830_ (.I0(\u_cpu.rf_ram.memory[8][7] ),
    .I1(\u_cpu.rf_ram.memory[9][7] ),
    .I2(\u_cpu.rf_ram.memory[10][7] ),
    .I3(\u_cpu.rf_ram.memory[11][7] ),
    .S0(_01591_),
    .S1(_01592_),
    .Z(_02440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06831_ (.A1(_01637_),
    .A2(_02440_),
    .ZN(_02441_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06832_ (.I0(\u_cpu.rf_ram.memory[12][7] ),
    .I1(\u_cpu.rf_ram.memory[13][7] ),
    .I2(\u_cpu.rf_ram.memory[14][7] ),
    .I3(\u_cpu.rf_ram.memory[15][7] ),
    .S0(_01813_),
    .S1(_01815_),
    .Z(_02442_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06833_ (.A1(_01399_),
    .A2(_02442_),
    .B(_02069_),
    .ZN(_02443_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06834_ (.I0(\u_cpu.rf_ram.memory[4][7] ),
    .I1(\u_cpu.rf_ram.memory[5][7] ),
    .I2(\u_cpu.rf_ram.memory[6][7] ),
    .I3(\u_cpu.rf_ram.memory[7][7] ),
    .S0(_01640_),
    .S1(_02071_),
    .Z(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06835_ (.A1(_01580_),
    .A2(_02444_),
    .ZN(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06836_ (.I0(\u_cpu.rf_ram.memory[0][7] ),
    .I1(\u_cpu.rf_ram.memory[1][7] ),
    .I2(\u_cpu.rf_ram.memory[2][7] ),
    .I3(\u_cpu.rf_ram.memory[3][7] ),
    .S0(_02074_),
    .S1(_01585_),
    .Z(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06837_ (.A1(_01786_),
    .A2(_02446_),
    .B(_01795_),
    .ZN(_02447_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06838_ (.A1(_02441_),
    .A2(_02443_),
    .B1(_02445_),
    .B2(_02447_),
    .C(_01807_),
    .ZN(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06839_ (.I0(\u_cpu.rf_ram.memory[20][7] ),
    .I1(\u_cpu.rf_ram.memory[21][7] ),
    .I2(\u_cpu.rf_ram.memory[22][7] ),
    .I3(\u_cpu.rf_ram.memory[23][7] ),
    .S0(_01631_),
    .S1(_01634_),
    .Z(_02449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06840_ (.A1(_02078_),
    .A2(_02449_),
    .ZN(_02450_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06841_ (.I0(\u_cpu.rf_ram.memory[16][7] ),
    .I1(\u_cpu.rf_ram.memory[17][7] ),
    .I2(\u_cpu.rf_ram.memory[18][7] ),
    .I3(\u_cpu.rf_ram.memory[19][7] ),
    .S0(_01598_),
    .S1(_01599_),
    .Z(_02451_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06842_ (.A1(_02081_),
    .A2(_02451_),
    .B(_01603_),
    .ZN(_02452_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06843_ (.I0(\u_cpu.rf_ram.memory[28][7] ),
    .I1(\u_cpu.rf_ram.memory[29][7] ),
    .I2(\u_cpu.rf_ram.memory[30][7] ),
    .I3(\u_cpu.rf_ram.memory[31][7] ),
    .S0(_02084_),
    .S1(_01577_),
    .Z(_02453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06844_ (.A1(_01590_),
    .A2(_02453_),
    .ZN(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06845_ (.I0(\u_cpu.rf_ram.memory[24][7] ),
    .I1(\u_cpu.rf_ram.memory[25][7] ),
    .I2(\u_cpu.rf_ram.memory[26][7] ),
    .I3(\u_cpu.rf_ram.memory[27][7] ),
    .S0(_01622_),
    .S1(_01625_),
    .Z(_02455_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06846_ (.A1(_01619_),
    .A2(_02455_),
    .B(_01588_),
    .ZN(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06847_ (.A1(_02450_),
    .A2(_02452_),
    .B1(_02454_),
    .B2(_02456_),
    .C(_01784_),
    .ZN(_02457_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06848_ (.I0(\u_cpu.rf_ram.memory[52][7] ),
    .I1(\u_cpu.rf_ram.memory[53][7] ),
    .I2(\u_cpu.rf_ram.memory[54][7] ),
    .I3(\u_cpu.rf_ram.memory[55][7] ),
    .S0(_01747_),
    .S1(_01748_),
    .Z(_02458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06849_ (.A1(_01697_),
    .A2(_02458_),
    .ZN(_02459_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06850_ (.I0(\u_cpu.rf_ram.memory[48][7] ),
    .I1(\u_cpu.rf_ram.memory[49][7] ),
    .I2(\u_cpu.rf_ram.memory[50][7] ),
    .I3(\u_cpu.rf_ram.memory[51][7] ),
    .S0(_01812_),
    .S1(_02092_),
    .Z(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06851_ (.A1(_01569_),
    .A2(_02460_),
    .B(_01602_),
    .ZN(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06852_ (.I0(\u_cpu.rf_ram.memory[60][7] ),
    .I1(\u_cpu.rf_ram.memory[61][7] ),
    .I2(\u_cpu.rf_ram.memory[62][7] ),
    .I3(\u_cpu.rf_ram.memory[63][7] ),
    .S0(_02095_),
    .S1(_01633_),
    .Z(_02462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06853_ (.A1(_01725_),
    .A2(_02462_),
    .ZN(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06854_ (.I0(\u_cpu.rf_ram.memory[56][7] ),
    .I1(\u_cpu.rf_ram.memory[57][7] ),
    .I2(\u_cpu.rf_ram.memory[58][7] ),
    .I3(\u_cpu.rf_ram.memory[59][7] ),
    .S0(_01729_),
    .S1(_02099_),
    .Z(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06855_ (.A1(_02098_),
    .A2(_02464_),
    .B(_01695_),
    .ZN(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06856_ (.A1(_02459_),
    .A2(_02461_),
    .B1(_02463_),
    .B2(_02465_),
    .C(_01427_),
    .ZN(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06857_ (.I0(\u_cpu.rf_ram.memory[40][7] ),
    .I1(\u_cpu.rf_ram.memory[41][7] ),
    .I2(\u_cpu.rf_ram.memory[42][7] ),
    .I3(\u_cpu.rf_ram.memory[43][7] ),
    .S0(_01736_),
    .S1(_02103_),
    .Z(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06858_ (.A1(_01772_),
    .A2(_02467_),
    .ZN(_02468_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06859_ (.I0(\u_cpu.rf_ram.memory[44][7] ),
    .I1(\u_cpu.rf_ram.memory[45][7] ),
    .I2(\u_cpu.rf_ram.memory[46][7] ),
    .I3(\u_cpu.rf_ram.memory[47][7] ),
    .S0(_01721_),
    .S1(_01624_),
    .Z(_02469_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06860_ (.A1(_01610_),
    .A2(_02469_),
    .B(_02107_),
    .ZN(_02470_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06861_ (.I0(\u_cpu.rf_ram.memory[36][7] ),
    .I1(\u_cpu.rf_ram.memory[37][7] ),
    .I2(\u_cpu.rf_ram.memory[38][7] ),
    .I3(\u_cpu.rf_ram.memory[39][7] ),
    .S0(_01716_),
    .S1(_02109_),
    .Z(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06862_ (.A1(_01715_),
    .A2(_02471_),
    .ZN(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06863_ (.I0(\u_cpu.rf_ram.memory[32][7] ),
    .I1(\u_cpu.rf_ram.memory[33][7] ),
    .I2(\u_cpu.rf_ram.memory[34][7] ),
    .I3(\u_cpu.rf_ram.memory[35][7] ),
    .S0(_01767_),
    .S1(_01768_),
    .Z(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06864_ (.A1(_01766_),
    .A2(_02473_),
    .B(_01731_),
    .ZN(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06865_ (.A1(_02468_),
    .A2(_02470_),
    .B1(_02472_),
    .B2(_02474_),
    .C(_01733_),
    .ZN(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06866_ (.A1(_01422_),
    .A2(_02466_),
    .A3(_02475_),
    .Z(_02476_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06867_ (.A1(_01760_),
    .A2(_02448_),
    .A3(_02457_),
    .B(_02476_),
    .ZN(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06868_ (.I0(\u_cpu.rf_ram.memory[108][7] ),
    .I1(\u_cpu.rf_ram.memory[109][7] ),
    .I2(\u_cpu.rf_ram.memory[110][7] ),
    .I3(\u_cpu.rf_ram.memory[111][7] ),
    .S0(_01639_),
    .S1(_01615_),
    .Z(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06869_ (.A1(_02117_),
    .A2(_02478_),
    .ZN(_02479_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06870_ (.I0(\u_cpu.rf_ram.memory[104][7] ),
    .I1(\u_cpu.rf_ram.memory[105][7] ),
    .I2(\u_cpu.rf_ram.memory[106][7] ),
    .I3(\u_cpu.rf_ram.memory[107][7] ),
    .S0(_01657_),
    .S1(_01660_),
    .Z(_02480_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06871_ (.A1(_01656_),
    .A2(_02480_),
    .B(_01587_),
    .ZN(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06872_ (.I0(\u_cpu.rf_ram.memory[100][7] ),
    .I1(\u_cpu.rf_ram.memory[101][7] ),
    .I2(\u_cpu.rf_ram.memory[102][7] ),
    .I3(\u_cpu.rf_ram.memory[103][7] ),
    .S0(_02122_),
    .S1(_01576_),
    .Z(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06873_ (.A1(_01802_),
    .A2(_02482_),
    .ZN(_02483_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06874_ (.I0(\u_cpu.rf_ram.memory[96][7] ),
    .I1(\u_cpu.rf_ram.memory[97][7] ),
    .I2(\u_cpu.rf_ram.memory[98][7] ),
    .I3(\u_cpu.rf_ram.memory[99][7] ),
    .S0(_02125_),
    .S1(_01693_),
    .Z(_02484_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06875_ (.A1(_01720_),
    .A2(_02484_),
    .B(_01663_),
    .ZN(_02485_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06876_ (.A1(_02479_),
    .A2(_02481_),
    .B1(_02483_),
    .B2(_02485_),
    .C(_01606_),
    .ZN(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06877_ (.I0(\u_cpu.rf_ram.memory[124][7] ),
    .I1(\u_cpu.rf_ram.memory[125][7] ),
    .I2(\u_cpu.rf_ram.memory[126][7] ),
    .I3(\u_cpu.rf_ram.memory[127][7] ),
    .S0(_01773_),
    .S1(_01774_),
    .Z(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06878_ (.A1(_01649_),
    .A2(_02487_),
    .ZN(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06879_ (.I0(\u_cpu.rf_ram.memory[120][7] ),
    .I1(\u_cpu.rf_ram.memory[121][7] ),
    .I2(\u_cpu.rf_ram.memory[122][7] ),
    .I3(\u_cpu.rf_ram.memory[123][7] ),
    .S0(_01674_),
    .S1(_01676_),
    .Z(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06880_ (.A1(_01672_),
    .A2(_02489_),
    .B(_01679_),
    .ZN(_02490_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06881_ (.I0(\u_cpu.rf_ram.memory[112][7] ),
    .I1(\u_cpu.rf_ram.memory[113][7] ),
    .I2(\u_cpu.rf_ram.memory[114][7] ),
    .I3(\u_cpu.rf_ram.memory[115][7] ),
    .S0(_02133_),
    .S1(_01699_),
    .Z(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06882_ (.A1(_01703_),
    .A2(_02491_),
    .ZN(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06883_ (.I0(\u_cpu.rf_ram.memory[116][7] ),
    .I1(\u_cpu.rf_ram.memory[117][7] ),
    .I2(\u_cpu.rf_ram.memory[118][7] ),
    .I3(\u_cpu.rf_ram.memory[119][7] ),
    .S0(_02136_),
    .S1(_01707_),
    .Z(_02493_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06884_ (.A1(_01691_),
    .A2(_02493_),
    .B(_01709_),
    .ZN(_02494_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06885_ (.A1(_02488_),
    .A2(_02490_),
    .B1(_02492_),
    .B2(_02494_),
    .C(_02139_),
    .ZN(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06886_ (.A1(_01647_),
    .A2(_02486_),
    .A3(_02495_),
    .ZN(_02496_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06887_ (.I0(\u_cpu.rf_ram.memory[92][7] ),
    .I1(\u_cpu.rf_ram.memory[93][7] ),
    .I2(\u_cpu.rf_ram.memory[94][7] ),
    .I3(\u_cpu.rf_ram.memory[95][7] ),
    .S0(_02142_),
    .S1(_01688_),
    .Z(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06888_ (.A1(_01735_),
    .A2(_02497_),
    .ZN(_02498_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06889_ (.I0(\u_cpu.rf_ram.memory[88][7] ),
    .I1(\u_cpu.rf_ram.memory[89][7] ),
    .I2(\u_cpu.rf_ram.memory[90][7] ),
    .I3(\u_cpu.rf_ram.memory[91][7] ),
    .S0(_01741_),
    .S1(_01742_),
    .Z(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06890_ (.A1(_01740_),
    .A2(_02499_),
    .B(_01744_),
    .ZN(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06891_ (.I0(\u_cpu.rf_ram.memory[80][7] ),
    .I1(\u_cpu.rf_ram.memory[81][7] ),
    .I2(\u_cpu.rf_ram.memory[82][7] ),
    .I3(\u_cpu.rf_ram.memory[83][7] ),
    .S0(_01651_),
    .S1(_01653_),
    .Z(_02501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06892_ (.A1(_02147_),
    .A2(_02501_),
    .ZN(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06893_ (.I0(\u_cpu.rf_ram.memory[84][7] ),
    .I1(\u_cpu.rf_ram.memory[85][7] ),
    .I2(\u_cpu.rf_ram.memory[86][7] ),
    .I3(\u_cpu.rf_ram.memory[87][7] ),
    .S0(_01752_),
    .S1(_02151_),
    .Z(_02503_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06894_ (.A1(_02150_),
    .A2(_02503_),
    .B(_02153_),
    .ZN(_02504_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06895_ (.A1(_02498_),
    .A2(_02500_),
    .B1(_02502_),
    .B2(_02504_),
    .C(_01757_),
    .ZN(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06896_ (.I0(\u_cpu.rf_ram.memory[64][7] ),
    .I1(\u_cpu.rf_ram.memory[65][7] ),
    .I2(\u_cpu.rf_ram.memory[66][7] ),
    .I3(\u_cpu.rf_ram.memory[67][7] ),
    .S0(_01798_),
    .S1(_01799_),
    .Z(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06897_ (.A1(_01797_),
    .A2(_02506_),
    .ZN(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06898_ (.I0(\u_cpu.rf_ram.memory[68][7] ),
    .I1(\u_cpu.rf_ram.memory[69][7] ),
    .I2(\u_cpu.rf_ram.memory[70][7] ),
    .I3(\u_cpu.rf_ram.memory[71][7] ),
    .S0(_01779_),
    .S1(_01780_),
    .Z(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06899_ (.A1(_01778_),
    .A2(_02508_),
    .B(_01782_),
    .ZN(_02509_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06900_ (.I0(\u_cpu.rf_ram.memory[72][7] ),
    .I1(\u_cpu.rf_ram.memory[73][7] ),
    .I2(\u_cpu.rf_ram.memory[74][7] ),
    .I3(\u_cpu.rf_ram.memory[75][7] ),
    .S0(_01762_),
    .S1(_01763_),
    .Z(_02510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06901_ (.A1(_01684_),
    .A2(_02510_),
    .ZN(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06902_ (.I0(\u_cpu.rf_ram.memory[76][7] ),
    .I1(\u_cpu.rf_ram.memory[77][7] ),
    .I2(\u_cpu.rf_ram.memory[78][7] ),
    .I3(\u_cpu.rf_ram.memory[79][7] ),
    .S0(_01792_),
    .S1(_01793_),
    .Z(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06903_ (.A1(_01791_),
    .A2(_02512_),
    .B(_01770_),
    .ZN(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06904_ (.A1(_02507_),
    .A2(_02509_),
    .B1(_02511_),
    .B2(_02513_),
    .C(_01711_),
    .ZN(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06905_ (.A1(_01565_),
    .A2(_02505_),
    .A3(_02514_),
    .ZN(_02515_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06906_ (.A1(_02496_),
    .A2(_02515_),
    .B(_01404_),
    .ZN(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06907_ (.I0(\u_cpu.rf_ram.memory[136][7] ),
    .I1(\u_cpu.rf_ram.memory[137][7] ),
    .I2(\u_cpu.rf_ram.memory[138][7] ),
    .I3(\u_cpu.rf_ram.memory[139][7] ),
    .S0(_01831_),
    .S1(_01832_),
    .Z(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06908_ (.A1(_01825_),
    .A2(_02517_),
    .ZN(_02518_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06909_ (.I0(\u_cpu.rf_ram.memory[140][7] ),
    .I1(\u_cpu.rf_ram.memory[141][7] ),
    .I2(\u_cpu.rf_ram.memory[142][7] ),
    .I3(\u_cpu.rf_ram.memory[143][7] ),
    .S0(_02169_),
    .S1(_01816_),
    .Z(_02519_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06910_ (.A1(_01830_),
    .A2(_02519_),
    .B(_01628_),
    .ZN(_02520_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06911_ (.I0(\u_cpu.rf_ram.memory[128][7] ),
    .I1(\u_cpu.rf_ram.memory[129][7] ),
    .I2(\u_cpu.rf_ram.memory[130][7] ),
    .I3(\u_cpu.rf_ram.memory[131][7] ),
    .S0(_01614_),
    .S1(_01616_),
    .Z(_02521_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06912_ (.A1(_01611_),
    .A2(_02521_),
    .ZN(_02522_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06913_ (.I0(\u_cpu.rf_ram.memory[132][7] ),
    .I1(\u_cpu.rf_ram.memory[133][7] ),
    .I2(\u_cpu.rf_ram.memory[134][7] ),
    .I3(\u_cpu.rf_ram.memory[135][7] ),
    .S0(_01826_),
    .S1(_02174_),
    .Z(_02523_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06914_ (.A1(_01570_),
    .A2(_02523_),
    .B(_01644_),
    .ZN(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _06915_ (.A1(_02518_),
    .A2(_02520_),
    .B1(_02522_),
    .B2(_02524_),
    .C(_01405_),
    .ZN(_02525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06916_ (.A1(_02516_),
    .A2(_02525_),
    .ZN(_02526_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06917_ (.A1(_01406_),
    .A2(_02477_),
    .B(_02526_),
    .ZN(_00007_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _06918_ (.A1(\u_cpu.cpu.state.o_cnt_r[0] ),
    .A2(\u_cpu.cpu.state.o_cnt_r[1] ),
    .A3(\u_cpu.cpu.state.o_cnt_r[2] ),
    .A4(\u_cpu.cpu.state.o_cnt_r[3] ),
    .Z(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06919_ (.I(_02527_),
    .Z(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06920_ (.I(_02528_),
    .Z(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06921_ (.I(_02529_),
    .Z(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06922_ (.I(_01410_),
    .ZN(_02531_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06923_ (.I(\u_cpu.cpu.branch_op ),
    .Z(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06924_ (.A1(\u_arbiter.i_wb_cpu_dbus_we ),
    .A2(\u_cpu.cpu.bufreg.i_sh_signed ),
    .B(_02531_),
    .C(_02532_),
    .ZN(_02533_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06925_ (.A1(\u_cpu.cpu.alu.i_rs1 ),
    .A2(\u_cpu.cpu.alu.add_cy_r ),
    .ZN(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06926_ (.I(\u_cpu.cpu.immdec.imm11_7[0] ),
    .ZN(_02535_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06927_ (.A1(\u_cpu.cpu.decode.opcode[2] ),
    .A2(\u_cpu.cpu.decode.opcode[1] ),
    .A3(\u_cpu.cpu.decode.opcode[0] ),
    .ZN(_02536_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06928_ (.A1(\u_arbiter.i_wb_cpu_dbus_we ),
    .A2(_02535_),
    .A3(_02536_),
    .Z(_02537_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06929_ (.A1(\u_arbiter.i_wb_cpu_dbus_we ),
    .A2(_02536_),
    .B(\u_cpu.cpu.immdec.imm24_20[0] ),
    .ZN(_02538_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06930_ (.A1(\u_cpu.cpu.csr_d_sel ),
    .A2(\u_cpu.cpu.decode.opcode[2] ),
    .A3(\u_cpu.cpu.branch_op ),
    .ZN(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06931_ (.A1(\u_cpu.cpu.bufreg2.i_cnt_done ),
    .A2(\u_cpu.cpu.immdec.imm31 ),
    .A3(_02539_),
    .ZN(_02540_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06932_ (.A1(\u_cpu.cpu.bufreg2.i_cnt_done ),
    .A2(_02537_),
    .A3(_02538_),
    .B(_02540_),
    .ZN(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06933_ (.I(\u_cpu.rf_ram.regzero ),
    .ZN(_02542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06934_ (.A1(\u_cpu.rf_ram.rdata[0] ),
    .A2(_02542_),
    .ZN(_02543_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06935_ (.A1(\u_cpu.rf_ram_if.rdata1[0] ),
    .A2(\u_cpu.rf_ram_if.rtrig1 ),
    .ZN(_02544_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06936_ (.A1(\u_cpu.rf_ram_if.rtrig1 ),
    .A2(_02543_),
    .B(_02544_),
    .ZN(_02545_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06937_ (.I0(_02541_),
    .I1(_02545_),
    .S(\u_arbiter.i_wb_cpu_dbus_we ),
    .Z(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06938_ (.I(_02546_),
    .Z(_02547_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06939_ (.A1(_02533_),
    .A2(_02547_),
    .Z(_02548_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06940_ (.I(\u_cpu.cpu.alu.i_rs1 ),
    .Z(_02549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06941_ (.A1(_02549_),
    .A2(\u_cpu.cpu.alu.add_cy_r ),
    .ZN(_02550_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06942_ (.A1(_02534_),
    .A2(_02548_),
    .B(_02550_),
    .ZN(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06943_ (.A1(_02530_),
    .A2(_02551_),
    .ZN(_02552_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06944_ (.A1(_02530_),
    .A2(_02533_),
    .B(_02552_),
    .ZN(_00021_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06945_ (.I(_01408_),
    .Z(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06946_ (.A1(_02553_),
    .A2(_01391_),
    .ZN(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06947_ (.A1(_02553_),
    .A2(_02549_),
    .B(_02554_),
    .ZN(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06948_ (.I(_01371_),
    .ZN(_02556_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06949_ (.I(_01372_),
    .ZN(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06950_ (.A1(_02556_),
    .A2(_02557_),
    .ZN(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06951_ (.I(_01371_),
    .Z(_02559_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06952_ (.A1(_02559_),
    .A2(_02555_),
    .B(_02557_),
    .ZN(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06953_ (.A1(_01380_),
    .A2(_01383_),
    .Z(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06954_ (.I(\u_cpu.cpu.decode.op22 ),
    .ZN(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06955_ (.I(\u_cpu.cpu.state.o_cnt_r[3] ),
    .Z(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06956_ (.A1(\u_cpu.cpu.mem_bytecnt[1] ),
    .A2(\u_cpu.cpu.state.o_cnt[2] ),
    .A3(\u_cpu.cpu.mem_bytecnt[0] ),
    .ZN(_02564_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06957_ (.I(_02564_),
    .Z(_02565_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06958_ (.A1(\u_cpu.cpu.decode.op26 ),
    .A2(_01413_),
    .ZN(_02566_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _06959_ (.A1(_02562_),
    .A2(_02563_),
    .A3(_02565_),
    .A4(_02566_),
    .Z(_02567_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06960_ (.I(\u_cpu.cpu.genblk3.csr.mcause3_0[0] ),
    .ZN(_02568_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06961_ (.I(\u_cpu.cpu.bufreg2.i_cnt_done ),
    .Z(_02569_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06962_ (.A1(_02569_),
    .A2(\u_cpu.cpu.genblk3.csr.mcause31 ),
    .B(_02564_),
    .ZN(_02570_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06963_ (.I(\u_cpu.cpu.decode.op21 ),
    .ZN(_02571_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06964_ (.A1(_02571_),
    .A2(\u_cpu.cpu.decode.co_ebreak ),
    .A3(_01413_),
    .ZN(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06965_ (.A1(_02528_),
    .A2(_02572_),
    .ZN(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _06966_ (.A1(_02568_),
    .A2(_02565_),
    .B(_02570_),
    .C(_02573_),
    .ZN(_02574_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _06967_ (.A1(_02561_),
    .A2(_02545_),
    .B1(_02567_),
    .B2(\u_cpu.cpu.genblk3.csr.mstatus_mie ),
    .C(_02574_),
    .ZN(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _06968_ (.A1(_01411_),
    .A2(_02555_),
    .A3(_02558_),
    .B1(_02560_),
    .B2(_02575_),
    .ZN(_02576_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06969_ (.A1(_01394_),
    .A2(_02576_),
    .ZN(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06970_ (.I(_01387_),
    .Z(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06971_ (.I(_02578_),
    .Z(_02579_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06972_ (.A1(_01431_),
    .A2(_02579_),
    .ZN(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06973_ (.A1(_02577_),
    .A2(_02580_),
    .ZN(\u_cpu.cpu.o_wdata1 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06974_ (.A1(\u_cpu.cpu.alu.i_rs1 ),
    .A2(_02547_),
    .ZN(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06975_ (.A1(\u_cpu.cpu.alu.i_rs1 ),
    .A2(_02547_),
    .B(_01408_),
    .ZN(_02582_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06976_ (.A1(_01372_),
    .A2(_02581_),
    .B(_02582_),
    .ZN(_02583_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06977_ (.A1(_02559_),
    .A2(_02581_),
    .B(_02583_),
    .ZN(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06978_ (.I(\u_cpu.cpu.alu.cmp_r ),
    .ZN(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06979_ (.A1(\u_cpu.cpu.state.o_cnt_r[0] ),
    .A2(_02565_),
    .ZN(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06980_ (.A1(_02553_),
    .A2(_02585_),
    .A3(_02586_),
    .ZN(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06981_ (.A1(\u_cpu.cpu.alu.i_rs1 ),
    .A2(\u_cpu.cpu.alu.add_cy_r ),
    .Z(_02588_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06982_ (.A1(_02588_),
    .A2(_02533_),
    .A3(_02546_),
    .Z(_02589_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06983_ (.A1(_01412_),
    .A2(_02589_),
    .ZN(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06984_ (.I(_01369_),
    .ZN(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06985_ (.A1(_01385_),
    .A2(\u_cpu.cpu.state.init_done ),
    .A3(_01386_),
    .A4(_01376_),
    .ZN(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06986_ (.A1(\u_cpu.cpu.branch_op ),
    .A2(\u_cpu.cpu.decode.opcode[0] ),
    .Z(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06987_ (.A1(_01408_),
    .A2(_01371_),
    .Z(_02594_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06988_ (.A1(_01411_),
    .A2(_02593_),
    .A3(_02594_),
    .B(_01374_),
    .ZN(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06989_ (.A1(_02527_),
    .A2(_02592_),
    .A3(_02595_),
    .ZN(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06990_ (.I(\u_cpu.cpu.state.init_done ),
    .Z(_02597_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06991_ (.A1(_01375_),
    .A2(_01371_),
    .ZN(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06992_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .A2(_01408_),
    .ZN(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06993_ (.A1(\u_cpu.cpu.state.stage_two_req ),
    .A2(_02599_),
    .ZN(_02600_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06994_ (.A1(_02597_),
    .A2(_02598_),
    .A3(_02600_),
    .ZN(_02601_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06995_ (.A1(_02596_),
    .A2(_02601_),
    .Z(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06996_ (.A1(_02591_),
    .A2(_02602_),
    .ZN(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06997_ (.A1(_02559_),
    .A2(_02587_),
    .B(_02590_),
    .C(_02603_),
    .ZN(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06998_ (.I(_01375_),
    .Z(_02605_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06999_ (.A1(_02584_),
    .A2(_02604_),
    .B(_02605_),
    .C(_02593_),
    .ZN(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07000_ (.I(\u_cpu.cpu.state.o_cnt_r[1] ),
    .ZN(_02607_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07001_ (.A1(\u_cpu.cpu.state.o_cnt_r[2] ),
    .A2(\u_cpu.cpu.ctrl.i_iscomp ),
    .ZN(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07002_ (.A1(_02607_),
    .A2(\u_cpu.cpu.ctrl.i_iscomp ),
    .B(_02608_),
    .ZN(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07003_ (.A1(_02564_),
    .A2(_02609_),
    .Z(_02610_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07004_ (.A1(\u_arbiter.i_wb_cpu_ibus_adr[0] ),
    .A2(\u_cpu.cpu.ctrl.pc_plus_4_cy_r ),
    .Z(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07005_ (.A1(_02610_),
    .A2(_02611_),
    .ZN(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07006_ (.I(_02532_),
    .Z(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07007_ (.I(\u_cpu.cpu.decode.opcode[0] ),
    .Z(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07008_ (.A1(_02613_),
    .A2(_02614_),
    .ZN(_02615_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07009_ (.I(_02614_),
    .ZN(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07010_ (.I(\u_cpu.cpu.mem_if.signbit ),
    .ZN(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07011_ (.A1(_02556_),
    .A2(\u_cpu.cpu.mem_bytecnt[1] ),
    .B1(\u_cpu.cpu.mem_bytecnt[0] ),
    .B2(_01411_),
    .ZN(_02618_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07012_ (.I0(\u_arbiter.i_wb_cpu_dbus_dat[0] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[8] ),
    .I2(\u_arbiter.i_wb_cpu_dbus_dat[16] ),
    .I3(\u_arbiter.i_wb_cpu_dbus_dat[24] ),
    .S0(\u_cpu.cpu.bufreg.lsb[0] ),
    .S1(\u_cpu.cpu.bufreg.lsb[1] ),
    .Z(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07013_ (.A1(_02618_),
    .A2(_02619_),
    .ZN(_02620_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07014_ (.A1(_02617_),
    .A2(_02618_),
    .B(_02620_),
    .ZN(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07015_ (.A1(_02553_),
    .A2(_02620_),
    .ZN(_02621_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07016_ (.A1(_02605_),
    .A2(_02616_),
    .A3(_00728_),
    .A4(_02621_),
    .ZN(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07017_ (.A1(_02612_),
    .A2(_02615_),
    .B(_02575_),
    .C(_02622_),
    .ZN(_02623_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07018_ (.A1(_01374_),
    .A2(_02614_),
    .ZN(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07019_ (.A1(\u_cpu.cpu.immdec.imm31 ),
    .A2(_02539_),
    .Z(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07020_ (.A1(_02569_),
    .A2(_02537_),
    .A3(_02538_),
    .ZN(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07021_ (.A1(_02569_),
    .A2(_02625_),
    .B(_02626_),
    .ZN(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07022_ (.A1(\u_cpu.cpu.state.o_cnt[2] ),
    .A2(\u_cpu.cpu.mem_bytecnt[0] ),
    .Z(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07023_ (.A1(_02532_),
    .A2(_02624_),
    .ZN(_02629_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07024_ (.A1(\u_cpu.cpu.mem_bytecnt[1] ),
    .A2(_02628_),
    .B(_02629_),
    .ZN(_02630_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07025_ (.A1(_02627_),
    .A2(_02630_),
    .ZN(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07026_ (.A1(_02591_),
    .A2(_02629_),
    .A3(_02602_),
    .ZN(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07027_ (.I(\u_arbiter.i_wb_cpu_dbus_we ),
    .Z(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07028_ (.A1(\u_cpu.cpu.decode.opcode[1] ),
    .A2(\u_cpu.cpu.decode.opcode[0] ),
    .B(_02536_),
    .ZN(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _07029_ (.A1(_02532_),
    .A2(_02633_),
    .B1(_01382_),
    .B2(_01379_),
    .C(_02634_),
    .ZN(_02635_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07030_ (.A1(\u_arbiter.i_wb_cpu_ibus_adr[0] ),
    .A2(_02635_),
    .ZN(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07031_ (.A1(\u_cpu.cpu.ctrl.pc_plus_offset_cy_r ),
    .A2(_02636_),
    .ZN(_02637_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07032_ (.A1(_02631_),
    .A2(_02632_),
    .B(_02637_),
    .ZN(_02638_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _07033_ (.A1(_02637_),
    .A2(_02631_),
    .A3(_02632_),
    .Z(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07034_ (.A1(_02638_),
    .A2(_02586_),
    .A3(_02639_),
    .ZN(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07035_ (.A1(_02613_),
    .A2(_02624_),
    .A3(_02640_),
    .ZN(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07036_ (.A1(_02606_),
    .A2(_02623_),
    .A3(_02641_),
    .ZN(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07037_ (.A1(_02613_),
    .A2(_02640_),
    .ZN(_02643_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07038_ (.A1(_02613_),
    .A2(_02603_),
    .B(_02643_),
    .C(_02578_),
    .ZN(_02644_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07039_ (.A1(_02579_),
    .A2(_02642_),
    .B(_02644_),
    .ZN(_02645_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07040_ (.I(_02645_),
    .Z(\u_cpu.cpu.o_wdata0 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07041_ (.I(\u_cpu.rf_ram_if.rtrig1 ),
    .Z(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07042_ (.I(_02646_),
    .Z(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07043_ (.I(_02542_),
    .Z(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07044_ (.A1(_02648_),
    .A2(\u_cpu.rf_ram.rdata[1] ),
    .ZN(_02649_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07045_ (.I(_02646_),
    .Z(_02650_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07046_ (.A1(_02650_),
    .A2(\u_cpu.rf_ram_if.rdata1[1] ),
    .ZN(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07047_ (.A1(_02647_),
    .A2(_02649_),
    .B(_02651_),
    .ZN(_00015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07048_ (.A1(_02648_),
    .A2(\u_cpu.rf_ram.rdata[2] ),
    .ZN(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07049_ (.A1(_02650_),
    .A2(\u_cpu.rf_ram_if.rdata1[2] ),
    .ZN(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07050_ (.A1(_02647_),
    .A2(_02652_),
    .B(_02653_),
    .ZN(_00016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07051_ (.A1(_02648_),
    .A2(\u_cpu.rf_ram.rdata[3] ),
    .ZN(_02654_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07052_ (.A1(_02650_),
    .A2(\u_cpu.rf_ram_if.rdata1[3] ),
    .ZN(_02655_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07053_ (.A1(_02647_),
    .A2(_02654_),
    .B(_02655_),
    .ZN(_00017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07054_ (.A1(_02542_),
    .A2(\u_cpu.rf_ram.rdata[4] ),
    .ZN(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07055_ (.A1(_02646_),
    .A2(\u_cpu.rf_ram_if.rdata1[4] ),
    .ZN(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07056_ (.A1(_02647_),
    .A2(_02656_),
    .B(_02657_),
    .ZN(_00018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07057_ (.A1(_02542_),
    .A2(\u_cpu.rf_ram.rdata[5] ),
    .ZN(_02658_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07058_ (.A1(_02646_),
    .A2(\u_cpu.rf_ram_if.rdata1[5] ),
    .ZN(_02659_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07059_ (.A1(_02647_),
    .A2(_02658_),
    .B(_02659_),
    .ZN(_00019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07060_ (.A1(_02542_),
    .A2(\u_cpu.rf_ram.rdata[6] ),
    .ZN(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07061_ (.A1(_02646_),
    .A2(\u_cpu.rf_ram_if.rdata1[6] ),
    .ZN(_02661_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07062_ (.A1(_02650_),
    .A2(_02660_),
    .B(_02661_),
    .ZN(_00020_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07063_ (.I(_01401_),
    .Z(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07064_ (.A1(\u_cpu.rf_ram_if.rdata0[1] ),
    .A2(_02662_),
    .ZN(_02663_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07065_ (.A1(_01430_),
    .A2(_02543_),
    .B(_02663_),
    .ZN(_00008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07066_ (.A1(\u_cpu.rf_ram_if.rdata0[2] ),
    .A2(_02662_),
    .ZN(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07067_ (.A1(_01430_),
    .A2(_02649_),
    .B(_02664_),
    .ZN(_00009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07068_ (.I(_01401_),
    .Z(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07069_ (.A1(\u_cpu.rf_ram_if.rdata0[3] ),
    .A2(_02665_),
    .ZN(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07070_ (.A1(_01430_),
    .A2(_02652_),
    .B(_02666_),
    .ZN(_00010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07071_ (.A1(\u_cpu.rf_ram_if.rdata0[4] ),
    .A2(_02665_),
    .ZN(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07072_ (.A1(_01430_),
    .A2(_02654_),
    .B(_02667_),
    .ZN(_00011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07073_ (.A1(\u_cpu.rf_ram_if.rdata0[5] ),
    .A2(_02665_),
    .ZN(_02668_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07074_ (.A1(_02662_),
    .A2(_02656_),
    .B(_02668_),
    .ZN(_00012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07075_ (.A1(\u_cpu.rf_ram_if.rdata0[6] ),
    .A2(_02665_),
    .ZN(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07076_ (.A1(_02662_),
    .A2(_02658_),
    .B(_02669_),
    .ZN(_00013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07077_ (.A1(\u_cpu.rf_ram_if.rdata0[7] ),
    .A2(_02665_),
    .ZN(_02670_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07078_ (.A1(_02662_),
    .A2(_02660_),
    .B(_02670_),
    .ZN(_00014_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07079_ (.I(_02556_),
    .Z(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07080_ (.I(_01370_),
    .ZN(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07081_ (.A1(_02671_),
    .A2(_02672_),
    .B1(_01411_),
    .B2(_02591_),
    .ZN(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _07082_ (.A1(\u_cpu.cpu.state.o_cnt_r[0] ),
    .A2(\u_cpu.cpu.state.o_cnt_r[1] ),
    .A3(\u_cpu.cpu.state.o_cnt_r[2] ),
    .A4(_02563_),
    .ZN(_02674_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07083_ (.I(_01374_),
    .Z(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07084_ (.I(_02532_),
    .Z(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07085_ (.A1(_02675_),
    .A2(_02676_),
    .ZN(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07086_ (.A1(_02597_),
    .A2(_02674_),
    .A3(_02677_),
    .ZN(_02678_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07087_ (.A1(_02673_),
    .A2(_02678_),
    .B(_01456_),
    .ZN(\u_arbiter.o_wb_cpu_cyc ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07088_ (.I(_02633_),
    .ZN(_02679_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07089_ (.A1(_02679_),
    .A2(_01434_),
    .ZN(\u_arbiter.o_wb_cpu_we ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07090_ (.I(\u_cpu.cpu.decode.opcode[1] ),
    .Z(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07091_ (.A1(_02676_),
    .A2(_02680_),
    .ZN(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07092_ (.A1(_02613_),
    .A2(_02616_),
    .ZN(_02682_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07093_ (.A1(_02549_),
    .A2(\u_cpu.cpu.bufreg.c_r ),
    .A3(_02681_),
    .A4(_02682_),
    .ZN(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07094_ (.I(_01376_),
    .Z(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07095_ (.A1(_02680_),
    .A2(_02614_),
    .Z(_02685_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07096_ (.A1(_02684_),
    .A2(_02586_),
    .A3(_02685_),
    .ZN(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07097_ (.A1(_02549_),
    .A2(_02681_),
    .A3(_02682_),
    .ZN(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07098_ (.A1(\u_cpu.cpu.bufreg.c_r ),
    .A2(_02687_),
    .Z(_02688_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _07099_ (.A1(_02675_),
    .A2(_02627_),
    .A3(_02686_),
    .A4(_02688_),
    .Z(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07100_ (.I(_02602_),
    .Z(_02690_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07101_ (.I(_02690_),
    .Z(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07102_ (.A1(_02683_),
    .A2(_02689_),
    .B(_02691_),
    .ZN(_00022_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07103_ (.A1(_01431_),
    .A2(\u_cpu.cpu.ctrl.pc_plus_offset_cy_r ),
    .A3(_02635_),
    .ZN(_02692_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07104_ (.I(\u_cpu.cpu.genblk3.csr.o_new_irq ),
    .Z(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07105_ (.A1(_02693_),
    .A2(_02597_),
    .ZN(_02694_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07106_ (.A1(_02694_),
    .A2(_02595_),
    .ZN(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07107_ (.A1(_02528_),
    .A2(_02695_),
    .ZN(_02696_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07108_ (.A1(_02692_),
    .A2(_02638_),
    .B(_02696_),
    .ZN(_00024_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07109_ (.A1(_01431_),
    .A2(\u_cpu.cpu.ctrl.pc_plus_4_cy_r ),
    .ZN(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07110_ (.A1(_02610_),
    .A2(_02611_),
    .ZN(_02698_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07111_ (.A1(_02697_),
    .A2(_02698_),
    .B(_02696_),
    .ZN(_00023_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07112_ (.I(_02674_),
    .Z(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07113_ (.A1(_01388_),
    .A2(_02699_),
    .ZN(\u_cpu.cpu.o_wen1 ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07114_ (.I(\u_cpu.cpu.immdec.imm11_7[2] ),
    .Z(_02700_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07115_ (.I(\u_cpu.cpu.immdec.imm11_7[3] ),
    .Z(_02701_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _07116_ (.A1(\u_cpu.cpu.immdec.imm11_7[1] ),
    .A2(_02700_),
    .A3(_02701_),
    .A4(\u_cpu.cpu.immdec.imm11_7[0] ),
    .Z(_02702_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07117_ (.I(_02614_),
    .Z(_02703_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07118_ (.A1(_02633_),
    .A2(_02703_),
    .B(_02615_),
    .C(_02605_),
    .ZN(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07119_ (.I(_02695_),
    .Z(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07120_ (.A1(\u_cpu.cpu.immdec.imm11_7[4] ),
    .A2(_02702_),
    .B(_02704_),
    .C(_02705_),
    .ZN(_02706_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07121_ (.A1(_01394_),
    .A2(_02706_),
    .B(_02699_),
    .ZN(\u_cpu.cpu.o_wen0 ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07122_ (.A1(_01369_),
    .A2(_01372_),
    .ZN(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07123_ (.A1(_01370_),
    .A2(_02707_),
    .B(_02671_),
    .ZN(\u_arbiter.i_wb_cpu_dbus_sel[1] ));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07124_ (.A1(_01369_),
    .A2(_02672_),
    .B(_02671_),
    .ZN(\u_arbiter.i_wb_cpu_dbus_sel[2] ));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07125_ (.A1(_02672_),
    .A2(_02707_),
    .B(_02671_),
    .ZN(\u_arbiter.i_wb_cpu_dbus_sel[3] ));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07126_ (.A1(_01387_),
    .A2(_01395_),
    .B(\u_cpu.rf_ram_if.genblk1.wtrig0_r ),
    .ZN(_02708_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07127_ (.A1(\u_cpu.rf_ram_if.genblk1.wtrig0_r ),
    .A2(_01387_),
    .ZN(_02709_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07128_ (.A1(_02535_),
    .A2(_02709_),
    .ZN(_02710_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07129_ (.A1(_02708_),
    .A2(_02710_),
    .ZN(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07130_ (.I(\u_cpu.rf_ram_if.genblk1.wtrig0_r ),
    .ZN(_02712_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07131_ (.A1(\u_cpu.cpu.immdec.imm11_7[1] ),
    .A2(_02712_),
    .ZN(_02713_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07132_ (.A1(_02712_),
    .A2(_01414_),
    .B(_02713_),
    .ZN(_02714_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07133_ (.A1(_02578_),
    .A2(_02714_),
    .ZN(_02715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07134_ (.A1(_02711_),
    .A2(_02715_),
    .ZN(_02716_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07135_ (.I(\u_cpu.rf_ram_if.rcnt[0] ),
    .Z(_02717_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07136_ (.A1(\u_cpu.rf_ram_if.rcnt[1] ),
    .A2(_02717_),
    .B(\u_cpu.rf_ram_if.rcnt[2] ),
    .ZN(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07137_ (.A1(\u_cpu.raddr[0] ),
    .A2(_02718_),
    .Z(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07138_ (.I(_02719_),
    .ZN(_02720_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07139_ (.A1(_01658_),
    .A2(_02720_),
    .ZN(_02721_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07140_ (.A1(_02716_),
    .A2(_02721_),
    .ZN(_02722_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07141_ (.I(_02722_),
    .Z(_02723_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07142_ (.I(_02709_),
    .Z(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07143_ (.A1(\u_cpu.cpu.immdec.imm11_7[2] ),
    .A2(_02724_),
    .ZN(_02725_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07144_ (.I(\u_cpu.rf_ram_if.genblk1.wtrig0_r ),
    .Z(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07145_ (.A1(_02726_),
    .A2(\u_cpu.rf_ram_if.wen1_r ),
    .B1(\u_cpu.rf_ram_if.rtrig0 ),
    .B2(\u_cpu.rf_ram_if.wen0_r ),
    .ZN(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07146_ (.I(_02727_),
    .ZN(_02728_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07147_ (.A1(\u_cpu.cpu.immdec.imm11_7[4] ),
    .A2(_02724_),
    .A3(_02728_),
    .ZN(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07148_ (.A1(_02701_),
    .A2(_02725_),
    .A3(_02729_),
    .ZN(_02730_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07149_ (.I(_02730_),
    .Z(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07150_ (.A1(_02723_),
    .A2(_02731_),
    .ZN(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07151_ (.I(_02732_),
    .Z(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07152_ (.I(_02712_),
    .Z(_02734_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07153_ (.I(_02734_),
    .Z(_02735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07154_ (.I(_02726_),
    .Z(_02736_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07155_ (.A1(\u_cpu.rf_ram_if.wdata1_r[0] ),
    .A2(_02736_),
    .Z(_02737_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07156_ (.A1(\u_cpu.rf_ram_if.wdata0_r[0] ),
    .A2(_02735_),
    .B(_02737_),
    .ZN(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07157_ (.I(_02738_),
    .Z(_02739_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07158_ (.I(_02739_),
    .Z(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07159_ (.I(_02732_),
    .Z(_02741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07160_ (.A1(\u_cpu.rf_ram.memory[82][0] ),
    .A2(_02741_),
    .ZN(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07161_ (.A1(_02733_),
    .A2(_02740_),
    .B(_02742_),
    .ZN(_00026_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07162_ (.A1(_02736_),
    .A2(\u_cpu.rf_ram_if.wdata1_r[1] ),
    .Z(_02743_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07163_ (.A1(_02735_),
    .A2(\u_cpu.rf_ram_if.wdata0_r[1] ),
    .B(_02743_),
    .ZN(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07164_ (.I(_02744_),
    .Z(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07165_ (.I(_02745_),
    .Z(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07166_ (.A1(\u_cpu.rf_ram.memory[82][1] ),
    .A2(_02741_),
    .ZN(_02747_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07167_ (.A1(_02733_),
    .A2(_02746_),
    .B(_02747_),
    .ZN(_00027_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07168_ (.I(_02726_),
    .Z(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07169_ (.A1(_02748_),
    .A2(\u_cpu.rf_ram_if.wdata1_r[2] ),
    .Z(_02749_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07170_ (.A1(_02735_),
    .A2(\u_cpu.rf_ram_if.wdata0_r[2] ),
    .B(_02749_),
    .ZN(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07171_ (.I(_02750_),
    .Z(_02751_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07172_ (.I(_02751_),
    .Z(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07173_ (.I(_02732_),
    .Z(_02753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07174_ (.A1(\u_cpu.rf_ram.memory[82][2] ),
    .A2(_02753_),
    .ZN(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07175_ (.A1(_02733_),
    .A2(_02752_),
    .B(_02754_),
    .ZN(_00028_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07176_ (.A1(_02748_),
    .A2(\u_cpu.rf_ram_if.wdata1_r[3] ),
    .Z(_02755_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07177_ (.A1(_02735_),
    .A2(\u_cpu.rf_ram_if.wdata0_r[3] ),
    .B(_02755_),
    .ZN(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07178_ (.I(_02756_),
    .Z(_02757_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07179_ (.I(_02757_),
    .Z(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07180_ (.A1(\u_cpu.rf_ram.memory[82][3] ),
    .A2(_02753_),
    .ZN(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07181_ (.A1(_02733_),
    .A2(_02758_),
    .B(_02759_),
    .ZN(_00029_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07182_ (.A1(_02748_),
    .A2(\u_cpu.rf_ram_if.wdata1_r[4] ),
    .Z(_02760_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07183_ (.A1(_02735_),
    .A2(\u_cpu.rf_ram_if.wdata0_r[4] ),
    .B(_02760_),
    .ZN(_02761_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07184_ (.I(_02761_),
    .Z(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07185_ (.I(_02762_),
    .Z(_02763_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07186_ (.A1(\u_cpu.rf_ram.memory[82][4] ),
    .A2(_02753_),
    .ZN(_02764_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07187_ (.A1(_02733_),
    .A2(_02763_),
    .B(_02764_),
    .ZN(_00030_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07188_ (.A1(_02748_),
    .A2(\u_cpu.rf_ram_if.wdata1_r[5] ),
    .Z(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07189_ (.A1(_02734_),
    .A2(\u_cpu.rf_ram_if.wdata0_r[5] ),
    .B(_02765_),
    .ZN(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07190_ (.I(_02766_),
    .Z(_02767_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07191_ (.I(_02767_),
    .Z(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07192_ (.A1(\u_cpu.rf_ram.memory[82][5] ),
    .A2(_02753_),
    .ZN(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07193_ (.A1(_02741_),
    .A2(_02768_),
    .B(_02769_),
    .ZN(_00031_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07194_ (.A1(_02748_),
    .A2(\u_cpu.rf_ram_if.wdata1_r[6] ),
    .Z(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07195_ (.A1(_02734_),
    .A2(\u_cpu.rf_ram_if.wdata0_r[6] ),
    .B(_02770_),
    .ZN(_02771_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07196_ (.I(_02771_),
    .Z(_02772_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07197_ (.I(_02772_),
    .Z(_02773_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07198_ (.A1(\u_cpu.rf_ram.memory[82][6] ),
    .A2(_02753_),
    .ZN(_02774_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07199_ (.A1(_02741_),
    .A2(_02773_),
    .B(_02774_),
    .ZN(_00032_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07200_ (.A1(_02726_),
    .A2(\u_cpu.rf_ram_if.wdata1_r[7] ),
    .Z(_02775_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07201_ (.A1(_02734_),
    .A2(\u_cpu.cpu.o_wdata0 ),
    .B(_02775_),
    .ZN(_02776_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07202_ (.I(_02776_),
    .Z(_02777_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07203_ (.I(_02777_),
    .Z(_02778_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07204_ (.A1(\u_cpu.rf_ram.memory[82][7] ),
    .A2(_02732_),
    .ZN(_02779_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07205_ (.A1(_02741_),
    .A2(_02778_),
    .B(_02779_),
    .ZN(_00033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07206_ (.A1(\u_cpu.rf_ram_if.rcnt[1] ),
    .A2(_02717_),
    .B(\u_cpu.raddr[0] ),
    .C(\u_cpu.rf_ram_if.rcnt[2] ),
    .ZN(_02780_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07207_ (.A1(\u_cpu.raddr[1] ),
    .A2(_02780_),
    .Z(_02781_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _07208_ (.A1(_02720_),
    .A2(_02781_),
    .Z(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07209_ (.A1(_02708_),
    .A2(_02710_),
    .Z(_02783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07210_ (.A1(_02783_),
    .A2(_02715_),
    .ZN(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07211_ (.A1(_02782_),
    .A2(_02784_),
    .ZN(_02785_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07212_ (.I(_02785_),
    .Z(_02786_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07213_ (.I(\u_cpu.cpu.immdec.imm11_7[4] ),
    .ZN(_02787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07214_ (.A1(_02787_),
    .A2(_02728_),
    .ZN(_02788_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07215_ (.A1(_02701_),
    .A2(_02725_),
    .A3(_02788_),
    .ZN(_02789_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07216_ (.I(_02789_),
    .Z(_02790_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07217_ (.A1(_02786_),
    .A2(_02790_),
    .ZN(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07218_ (.I(_02791_),
    .Z(_02792_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07219_ (.I(_02791_),
    .Z(_02793_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07220_ (.A1(\u_cpu.rf_ram.memory[21][0] ),
    .A2(_02793_),
    .ZN(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07221_ (.A1(_02740_),
    .A2(_02792_),
    .B(_02794_),
    .ZN(_00034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07222_ (.A1(\u_cpu.rf_ram.memory[21][1] ),
    .A2(_02793_),
    .ZN(_02795_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07223_ (.A1(_02746_),
    .A2(_02792_),
    .B(_02795_),
    .ZN(_00035_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07224_ (.I(_02791_),
    .Z(_02796_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07225_ (.A1(\u_cpu.rf_ram.memory[21][2] ),
    .A2(_02796_),
    .ZN(_02797_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07226_ (.A1(_02752_),
    .A2(_02792_),
    .B(_02797_),
    .ZN(_00036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07227_ (.A1(\u_cpu.rf_ram.memory[21][3] ),
    .A2(_02796_),
    .ZN(_02798_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07228_ (.A1(_02758_),
    .A2(_02792_),
    .B(_02798_),
    .ZN(_00037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07229_ (.A1(\u_cpu.rf_ram.memory[21][4] ),
    .A2(_02796_),
    .ZN(_02799_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07230_ (.A1(_02763_),
    .A2(_02792_),
    .B(_02799_),
    .ZN(_00038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07231_ (.A1(\u_cpu.rf_ram.memory[21][5] ),
    .A2(_02796_),
    .ZN(_02800_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07232_ (.A1(_02768_),
    .A2(_02793_),
    .B(_02800_),
    .ZN(_00039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07233_ (.A1(\u_cpu.rf_ram.memory[21][6] ),
    .A2(_02796_),
    .ZN(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07234_ (.A1(_02773_),
    .A2(_02793_),
    .B(_02801_),
    .ZN(_00040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07235_ (.A1(\u_cpu.rf_ram.memory[21][7] ),
    .A2(_02791_),
    .ZN(_02802_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07236_ (.A1(_02778_),
    .A2(_02793_),
    .B(_02802_),
    .ZN(_00041_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07237_ (.A1(_02716_),
    .A2(_02782_),
    .ZN(_02803_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07238_ (.I(_02803_),
    .Z(_02804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07239_ (.A1(_02731_),
    .A2(_02804_),
    .ZN(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07240_ (.I(_02805_),
    .Z(_02806_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07241_ (.I(_02805_),
    .Z(_02807_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07242_ (.A1(\u_cpu.rf_ram.memory[81][0] ),
    .A2(_02807_),
    .ZN(_02808_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07243_ (.A1(_02740_),
    .A2(_02806_),
    .B(_02808_),
    .ZN(_00042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07244_ (.A1(\u_cpu.rf_ram.memory[81][1] ),
    .A2(_02807_),
    .ZN(_02809_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07245_ (.A1(_02746_),
    .A2(_02806_),
    .B(_02809_),
    .ZN(_00043_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07246_ (.I(_02805_),
    .Z(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07247_ (.A1(\u_cpu.rf_ram.memory[81][2] ),
    .A2(_02810_),
    .ZN(_02811_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07248_ (.A1(_02752_),
    .A2(_02806_),
    .B(_02811_),
    .ZN(_00044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07249_ (.A1(\u_cpu.rf_ram.memory[81][3] ),
    .A2(_02810_),
    .ZN(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07250_ (.A1(_02758_),
    .A2(_02806_),
    .B(_02812_),
    .ZN(_00045_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07251_ (.A1(\u_cpu.rf_ram.memory[81][4] ),
    .A2(_02810_),
    .ZN(_02813_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07252_ (.A1(_02763_),
    .A2(_02806_),
    .B(_02813_),
    .ZN(_00046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07253_ (.A1(\u_cpu.rf_ram.memory[81][5] ),
    .A2(_02810_),
    .ZN(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07254_ (.A1(_02768_),
    .A2(_02807_),
    .B(_02814_),
    .ZN(_00047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07255_ (.A1(\u_cpu.rf_ram.memory[81][6] ),
    .A2(_02810_),
    .ZN(_02815_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07256_ (.A1(_02773_),
    .A2(_02807_),
    .B(_02815_),
    .ZN(_00048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07257_ (.A1(\u_cpu.rf_ram.memory[81][7] ),
    .A2(_02805_),
    .ZN(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07258_ (.A1(_02778_),
    .A2(_02807_),
    .B(_02816_),
    .ZN(_00049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07259_ (.A1(_02723_),
    .A2(_02790_),
    .ZN(_02817_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07260_ (.I(_02817_),
    .Z(_02818_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07261_ (.I(_02817_),
    .Z(_02819_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07262_ (.A1(\u_cpu.rf_ram.memory[18][0] ),
    .A2(_02819_),
    .ZN(_02820_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07263_ (.A1(_02740_),
    .A2(_02818_),
    .B(_02820_),
    .ZN(_00050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07264_ (.A1(\u_cpu.rf_ram.memory[18][1] ),
    .A2(_02819_),
    .ZN(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07265_ (.A1(_02746_),
    .A2(_02818_),
    .B(_02821_),
    .ZN(_00051_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07266_ (.I(_02817_),
    .Z(_02822_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07267_ (.A1(\u_cpu.rf_ram.memory[18][2] ),
    .A2(_02822_),
    .ZN(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07268_ (.A1(_02752_),
    .A2(_02818_),
    .B(_02823_),
    .ZN(_00052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07269_ (.A1(\u_cpu.rf_ram.memory[18][3] ),
    .A2(_02822_),
    .ZN(_02824_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07270_ (.A1(_02758_),
    .A2(_02818_),
    .B(_02824_),
    .ZN(_00053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07271_ (.A1(\u_cpu.rf_ram.memory[18][4] ),
    .A2(_02822_),
    .ZN(_02825_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07272_ (.A1(_02763_),
    .A2(_02818_),
    .B(_02825_),
    .ZN(_00054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07273_ (.A1(\u_cpu.rf_ram.memory[18][5] ),
    .A2(_02822_),
    .ZN(_02826_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07274_ (.A1(_02768_),
    .A2(_02819_),
    .B(_02826_),
    .ZN(_00055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07275_ (.A1(\u_cpu.rf_ram.memory[18][6] ),
    .A2(_02822_),
    .ZN(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07276_ (.A1(_02773_),
    .A2(_02819_),
    .B(_02827_),
    .ZN(_00056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07277_ (.A1(\u_cpu.rf_ram.memory[18][7] ),
    .A2(_02817_),
    .ZN(_02828_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07278_ (.A1(_02778_),
    .A2(_02819_),
    .B(_02828_),
    .ZN(_00057_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _07279_ (.A1(_01658_),
    .A2(_02719_),
    .Z(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07280_ (.A1(_02784_),
    .A2(_02829_),
    .ZN(_02830_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07281_ (.I(_02830_),
    .Z(_02831_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07282_ (.A1(_02790_),
    .A2(_02831_),
    .ZN(_02832_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07283_ (.I(_02832_),
    .Z(_02833_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07284_ (.I(_02832_),
    .Z(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07285_ (.A1(\u_cpu.rf_ram.memory[20][0] ),
    .A2(_02834_),
    .ZN(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07286_ (.A1(_02740_),
    .A2(_02833_),
    .B(_02835_),
    .ZN(_00058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07287_ (.A1(\u_cpu.rf_ram.memory[20][1] ),
    .A2(_02834_),
    .ZN(_02836_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07288_ (.A1(_02746_),
    .A2(_02833_),
    .B(_02836_),
    .ZN(_00059_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07289_ (.I(_02832_),
    .Z(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07290_ (.A1(\u_cpu.rf_ram.memory[20][2] ),
    .A2(_02837_),
    .ZN(_02838_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07291_ (.A1(_02752_),
    .A2(_02833_),
    .B(_02838_),
    .ZN(_00060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07292_ (.A1(\u_cpu.rf_ram.memory[20][3] ),
    .A2(_02837_),
    .ZN(_02839_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07293_ (.A1(_02758_),
    .A2(_02833_),
    .B(_02839_),
    .ZN(_00061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07294_ (.A1(\u_cpu.rf_ram.memory[20][4] ),
    .A2(_02837_),
    .ZN(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07295_ (.A1(_02763_),
    .A2(_02833_),
    .B(_02840_),
    .ZN(_00062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07296_ (.A1(\u_cpu.rf_ram.memory[20][5] ),
    .A2(_02837_),
    .ZN(_02841_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07297_ (.A1(_02768_),
    .A2(_02834_),
    .B(_02841_),
    .ZN(_00063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07298_ (.A1(\u_cpu.rf_ram.memory[20][6] ),
    .A2(_02837_),
    .ZN(_02842_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07299_ (.A1(_02773_),
    .A2(_02834_),
    .B(_02842_),
    .ZN(_00064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07300_ (.A1(\u_cpu.rf_ram.memory[20][7] ),
    .A2(_02832_),
    .ZN(_02843_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07301_ (.A1(_02778_),
    .A2(_02834_),
    .B(_02843_),
    .ZN(_00065_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07302_ (.I(_02736_),
    .Z(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07303_ (.I0(\u_cpu.rf_ram_if.wdata0_r[0] ),
    .I1(\u_cpu.rf_ram_if.wdata1_r[0] ),
    .S(_02844_),
    .Z(_02845_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07304_ (.I(_02845_),
    .Z(_02846_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07305_ (.A1(\u_cpu.cpu.immdec.imm11_7[3] ),
    .A2(_02724_),
    .ZN(_02847_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07306_ (.A1(_02725_),
    .A2(_02847_),
    .ZN(_02848_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _07307_ (.A1(_02726_),
    .A2(_02578_),
    .A3(_02788_),
    .A4(_02848_),
    .ZN(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07308_ (.I(_02849_),
    .Z(_02850_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07309_ (.A1(_02804_),
    .A2(_02850_),
    .ZN(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07310_ (.I(_02851_),
    .Z(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07311_ (.I0(_02846_),
    .I1(\u_cpu.rf_ram.memory[1][0] ),
    .S(_02852_),
    .Z(_02853_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07312_ (.I(_02853_),
    .Z(_00066_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07313_ (.I0(\u_cpu.rf_ram_if.wdata0_r[1] ),
    .I1(\u_cpu.rf_ram_if.wdata1_r[1] ),
    .S(_02844_),
    .Z(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07314_ (.I(_02854_),
    .Z(_02855_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07315_ (.I0(_02855_),
    .I1(\u_cpu.rf_ram.memory[1][1] ),
    .S(_02852_),
    .Z(_02856_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07316_ (.I(_02856_),
    .Z(_00067_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07317_ (.I0(\u_cpu.rf_ram_if.wdata0_r[2] ),
    .I1(\u_cpu.rf_ram_if.wdata1_r[2] ),
    .S(_02844_),
    .Z(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07318_ (.I(_02857_),
    .Z(_02858_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07319_ (.I0(_02858_),
    .I1(\u_cpu.rf_ram.memory[1][2] ),
    .S(_02852_),
    .Z(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07320_ (.I(_02859_),
    .Z(_00068_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07321_ (.I0(\u_cpu.rf_ram_if.wdata0_r[3] ),
    .I1(\u_cpu.rf_ram_if.wdata1_r[3] ),
    .S(_02844_),
    .Z(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07322_ (.I(_02860_),
    .Z(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07323_ (.I0(_02861_),
    .I1(\u_cpu.rf_ram.memory[1][3] ),
    .S(_02852_),
    .Z(_02862_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07324_ (.I(_02862_),
    .Z(_00069_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07325_ (.I0(\u_cpu.rf_ram_if.wdata0_r[4] ),
    .I1(\u_cpu.rf_ram_if.wdata1_r[4] ),
    .S(_02844_),
    .Z(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07326_ (.I(_02863_),
    .Z(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07327_ (.I0(_02864_),
    .I1(\u_cpu.rf_ram.memory[1][4] ),
    .S(_02852_),
    .Z(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07328_ (.I(_02865_),
    .Z(_00070_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07329_ (.I0(\u_cpu.rf_ram_if.wdata0_r[5] ),
    .I1(\u_cpu.rf_ram_if.wdata1_r[5] ),
    .S(_02736_),
    .Z(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07330_ (.I(_02866_),
    .Z(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07331_ (.I0(_02867_),
    .I1(\u_cpu.rf_ram.memory[1][5] ),
    .S(_02851_),
    .Z(_02868_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07332_ (.I(_02868_),
    .Z(_00071_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07333_ (.I0(\u_cpu.rf_ram_if.wdata0_r[6] ),
    .I1(\u_cpu.rf_ram_if.wdata1_r[6] ),
    .S(_02736_),
    .Z(_02869_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07334_ (.I(_02869_),
    .Z(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07335_ (.I0(_02870_),
    .I1(\u_cpu.rf_ram.memory[1][6] ),
    .S(_02851_),
    .Z(_02871_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07336_ (.I(_02871_),
    .Z(_00072_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07337_ (.I0(\u_cpu.rf_ram_if.wdata1_r[7] ),
    .I1(\u_cpu.cpu.o_wdata0 ),
    .S(_02734_),
    .Z(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07338_ (.I(_02872_),
    .Z(_02873_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07339_ (.I0(_02873_),
    .I1(\u_cpu.rf_ram.memory[1][7] ),
    .S(_02851_),
    .Z(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07340_ (.I(_02874_),
    .Z(_00073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07341_ (.A1(_02719_),
    .A2(_02781_),
    .ZN(_02875_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07342_ (.A1(_02784_),
    .A2(_02875_),
    .ZN(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07343_ (.I(_02876_),
    .Z(_02877_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07344_ (.A1(_02850_),
    .A2(_02877_),
    .ZN(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07345_ (.I(_02878_),
    .Z(_02879_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07346_ (.I0(_02846_),
    .I1(\u_cpu.rf_ram.memory[7][0] ),
    .S(_02879_),
    .Z(_02880_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07347_ (.I(_02880_),
    .Z(_00074_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07348_ (.I0(_02855_),
    .I1(\u_cpu.rf_ram.memory[7][1] ),
    .S(_02879_),
    .Z(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07349_ (.I(_02881_),
    .Z(_00075_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07350_ (.I0(_02858_),
    .I1(\u_cpu.rf_ram.memory[7][2] ),
    .S(_02879_),
    .Z(_02882_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07351_ (.I(_02882_),
    .Z(_00076_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07352_ (.I0(_02861_),
    .I1(\u_cpu.rf_ram.memory[7][3] ),
    .S(_02879_),
    .Z(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07353_ (.I(_02883_),
    .Z(_00077_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07354_ (.I0(_02864_),
    .I1(\u_cpu.rf_ram.memory[7][4] ),
    .S(_02879_),
    .Z(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07355_ (.I(_02884_),
    .Z(_00078_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07356_ (.I0(_02867_),
    .I1(\u_cpu.rf_ram.memory[7][5] ),
    .S(_02878_),
    .Z(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07357_ (.I(_02885_),
    .Z(_00079_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07358_ (.I0(_02870_),
    .I1(\u_cpu.rf_ram.memory[7][6] ),
    .S(_02878_),
    .Z(_02886_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07359_ (.I(_02886_),
    .Z(_00080_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07360_ (.I0(_02873_),
    .I1(\u_cpu.rf_ram.memory[7][7] ),
    .S(_02878_),
    .Z(_02887_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07361_ (.I(_02887_),
    .Z(_00081_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07362_ (.I(_02739_),
    .Z(_02888_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07363_ (.I(_02888_),
    .Z(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07364_ (.A1(_02716_),
    .A2(_02829_),
    .ZN(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07365_ (.I(_02890_),
    .Z(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07366_ (.A1(_02731_),
    .A2(_02891_),
    .ZN(_02892_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07367_ (.I(_02892_),
    .Z(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07368_ (.I(_02892_),
    .Z(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07369_ (.A1(\u_cpu.rf_ram.memory[80][0] ),
    .A2(_02894_),
    .ZN(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07370_ (.A1(_02889_),
    .A2(_02893_),
    .B(_02895_),
    .ZN(_00082_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07371_ (.I(_02745_),
    .Z(_02896_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07372_ (.I(_02896_),
    .Z(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07373_ (.A1(\u_cpu.rf_ram.memory[80][1] ),
    .A2(_02894_),
    .ZN(_02898_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07374_ (.A1(_02897_),
    .A2(_02893_),
    .B(_02898_),
    .ZN(_00083_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07375_ (.I(_02751_),
    .Z(_02899_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07376_ (.I(_02899_),
    .Z(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07377_ (.I(_02892_),
    .Z(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07378_ (.A1(\u_cpu.rf_ram.memory[80][2] ),
    .A2(_02901_),
    .ZN(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07379_ (.A1(_02900_),
    .A2(_02893_),
    .B(_02902_),
    .ZN(_00084_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07380_ (.I(_02757_),
    .Z(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07381_ (.I(_02903_),
    .Z(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07382_ (.A1(\u_cpu.rf_ram.memory[80][3] ),
    .A2(_02901_),
    .ZN(_02905_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07383_ (.A1(_02904_),
    .A2(_02893_),
    .B(_02905_),
    .ZN(_00085_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07384_ (.I(_02762_),
    .Z(_02906_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07385_ (.I(_02906_),
    .Z(_02907_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07386_ (.A1(\u_cpu.rf_ram.memory[80][4] ),
    .A2(_02901_),
    .ZN(_02908_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07387_ (.A1(_02907_),
    .A2(_02893_),
    .B(_02908_),
    .ZN(_00086_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07388_ (.I(_02767_),
    .Z(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07389_ (.I(_02909_),
    .Z(_02910_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07390_ (.A1(\u_cpu.rf_ram.memory[80][5] ),
    .A2(_02901_),
    .ZN(_02911_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07391_ (.A1(_02910_),
    .A2(_02894_),
    .B(_02911_),
    .ZN(_00087_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07392_ (.I(_02772_),
    .Z(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07393_ (.I(_02912_),
    .Z(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07394_ (.A1(\u_cpu.rf_ram.memory[80][6] ),
    .A2(_02901_),
    .ZN(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07395_ (.A1(_02913_),
    .A2(_02894_),
    .B(_02914_),
    .ZN(_00088_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07396_ (.I(_02777_),
    .Z(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07397_ (.I(_02915_),
    .Z(_02916_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07398_ (.A1(\u_cpu.rf_ram.memory[80][7] ),
    .A2(_02892_),
    .ZN(_02917_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07399_ (.A1(_02916_),
    .A2(_02894_),
    .B(_02917_),
    .ZN(_00089_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07400_ (.A1(_02578_),
    .A2(_02714_),
    .Z(_02918_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07401_ (.A1(_02783_),
    .A2(_02918_),
    .ZN(_02919_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07402_ (.A1(_02721_),
    .A2(_02919_),
    .ZN(_02920_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07403_ (.I(_02920_),
    .Z(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07404_ (.A1(_02729_),
    .A2(_02848_),
    .ZN(_02922_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07405_ (.I(_02922_),
    .Z(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07406_ (.A1(_02921_),
    .A2(_02923_),
    .ZN(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07407_ (.I(_02924_),
    .Z(_02925_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07408_ (.I(_02924_),
    .Z(_02926_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07409_ (.A1(\u_cpu.rf_ram.memory[78][0] ),
    .A2(_02926_),
    .ZN(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07410_ (.A1(_02889_),
    .A2(_02925_),
    .B(_02927_),
    .ZN(_00090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07411_ (.A1(\u_cpu.rf_ram.memory[78][1] ),
    .A2(_02926_),
    .ZN(_02928_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07412_ (.A1(_02897_),
    .A2(_02925_),
    .B(_02928_),
    .ZN(_00091_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07413_ (.I(_02924_),
    .Z(_02929_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07414_ (.A1(\u_cpu.rf_ram.memory[78][2] ),
    .A2(_02929_),
    .ZN(_02930_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07415_ (.A1(_02900_),
    .A2(_02925_),
    .B(_02930_),
    .ZN(_00092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07416_ (.A1(\u_cpu.rf_ram.memory[78][3] ),
    .A2(_02929_),
    .ZN(_02931_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07417_ (.A1(_02904_),
    .A2(_02925_),
    .B(_02931_),
    .ZN(_00093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07418_ (.A1(\u_cpu.rf_ram.memory[78][4] ),
    .A2(_02929_),
    .ZN(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07419_ (.A1(_02907_),
    .A2(_02925_),
    .B(_02932_),
    .ZN(_00094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07420_ (.A1(\u_cpu.rf_ram.memory[78][5] ),
    .A2(_02929_),
    .ZN(_02933_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07421_ (.A1(_02910_),
    .A2(_02926_),
    .B(_02933_),
    .ZN(_00095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07422_ (.A1(\u_cpu.rf_ram.memory[78][6] ),
    .A2(_02929_),
    .ZN(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07423_ (.A1(_02913_),
    .A2(_02926_),
    .B(_02934_),
    .ZN(_00096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07424_ (.A1(\u_cpu.rf_ram.memory[78][7] ),
    .A2(_02924_),
    .ZN(_02935_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07425_ (.A1(_02916_),
    .A2(_02926_),
    .B(_02935_),
    .ZN(_00097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07426_ (.A1(_02711_),
    .A2(_02918_),
    .ZN(_02936_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07427_ (.A1(_02721_),
    .A2(_02936_),
    .ZN(_02937_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07428_ (.I(_02937_),
    .Z(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07429_ (.A1(_02700_),
    .A2(_02788_),
    .A3(_02847_),
    .ZN(_02939_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07430_ (.I(_02939_),
    .Z(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07431_ (.A1(_02938_),
    .A2(_02940_),
    .ZN(_02941_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07432_ (.I(_02941_),
    .Z(_02942_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07433_ (.I(_02941_),
    .Z(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07434_ (.A1(\u_cpu.rf_ram.memory[42][0] ),
    .A2(_02943_),
    .ZN(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07435_ (.A1(_02889_),
    .A2(_02942_),
    .B(_02944_),
    .ZN(_00098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07436_ (.A1(\u_cpu.rf_ram.memory[42][1] ),
    .A2(_02943_),
    .ZN(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07437_ (.A1(_02897_),
    .A2(_02942_),
    .B(_02945_),
    .ZN(_00099_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07438_ (.I(_02941_),
    .Z(_02946_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07439_ (.A1(\u_cpu.rf_ram.memory[42][2] ),
    .A2(_02946_),
    .ZN(_02947_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07440_ (.A1(_02900_),
    .A2(_02942_),
    .B(_02947_),
    .ZN(_00100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07441_ (.A1(\u_cpu.rf_ram.memory[42][3] ),
    .A2(_02946_),
    .ZN(_02948_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07442_ (.A1(_02904_),
    .A2(_02942_),
    .B(_02948_),
    .ZN(_00101_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07443_ (.A1(\u_cpu.rf_ram.memory[42][4] ),
    .A2(_02946_),
    .ZN(_02949_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07444_ (.A1(_02907_),
    .A2(_02942_),
    .B(_02949_),
    .ZN(_00102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07445_ (.A1(\u_cpu.rf_ram.memory[42][5] ),
    .A2(_02946_),
    .ZN(_02950_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07446_ (.A1(_02910_),
    .A2(_02943_),
    .B(_02950_),
    .ZN(_00103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07447_ (.A1(\u_cpu.rf_ram.memory[42][6] ),
    .A2(_02946_),
    .ZN(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07448_ (.A1(_02913_),
    .A2(_02943_),
    .B(_02951_),
    .ZN(_00104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07449_ (.A1(\u_cpu.rf_ram.memory[42][7] ),
    .A2(_02941_),
    .ZN(_02952_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07450_ (.A1(_02916_),
    .A2(_02943_),
    .B(_02952_),
    .ZN(_00105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07451_ (.A1(_02921_),
    .A2(_02940_),
    .ZN(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07452_ (.I(_02953_),
    .Z(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07453_ (.I(_02953_),
    .Z(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07454_ (.A1(\u_cpu.rf_ram.memory[46][0] ),
    .A2(_02955_),
    .ZN(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07455_ (.A1(_02889_),
    .A2(_02954_),
    .B(_02956_),
    .ZN(_00106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07456_ (.A1(\u_cpu.rf_ram.memory[46][1] ),
    .A2(_02955_),
    .ZN(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07457_ (.A1(_02897_),
    .A2(_02954_),
    .B(_02957_),
    .ZN(_00107_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07458_ (.I(_02953_),
    .Z(_02958_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07459_ (.A1(\u_cpu.rf_ram.memory[46][2] ),
    .A2(_02958_),
    .ZN(_02959_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07460_ (.A1(_02900_),
    .A2(_02954_),
    .B(_02959_),
    .ZN(_00108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07461_ (.A1(\u_cpu.rf_ram.memory[46][3] ),
    .A2(_02958_),
    .ZN(_02960_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07462_ (.A1(_02904_),
    .A2(_02954_),
    .B(_02960_),
    .ZN(_00109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07463_ (.A1(\u_cpu.rf_ram.memory[46][4] ),
    .A2(_02958_),
    .ZN(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07464_ (.A1(_02907_),
    .A2(_02954_),
    .B(_02961_),
    .ZN(_00110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07465_ (.A1(\u_cpu.rf_ram.memory[46][5] ),
    .A2(_02958_),
    .ZN(_02962_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07466_ (.A1(_02910_),
    .A2(_02955_),
    .B(_02962_),
    .ZN(_00111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07467_ (.A1(\u_cpu.rf_ram.memory[46][6] ),
    .A2(_02958_),
    .ZN(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07468_ (.A1(_02913_),
    .A2(_02955_),
    .B(_02963_),
    .ZN(_00112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07469_ (.A1(\u_cpu.rf_ram.memory[46][7] ),
    .A2(_02953_),
    .ZN(_02964_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07470_ (.A1(_02916_),
    .A2(_02955_),
    .B(_02964_),
    .ZN(_00113_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07471_ (.I(_02939_),
    .Z(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07472_ (.A1(_02782_),
    .A2(_02919_),
    .ZN(_02966_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07473_ (.I(_02966_),
    .Z(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07474_ (.A1(_02965_),
    .A2(_02967_),
    .ZN(_02968_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07475_ (.I(_02968_),
    .Z(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07476_ (.I(_02968_),
    .Z(_02970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07477_ (.A1(\u_cpu.rf_ram.memory[45][0] ),
    .A2(_02970_),
    .ZN(_02971_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07478_ (.A1(_02889_),
    .A2(_02969_),
    .B(_02971_),
    .ZN(_00114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07479_ (.A1(\u_cpu.rf_ram.memory[45][1] ),
    .A2(_02970_),
    .ZN(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07480_ (.A1(_02897_),
    .A2(_02969_),
    .B(_02972_),
    .ZN(_00115_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07481_ (.I(_02968_),
    .Z(_02973_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07482_ (.A1(\u_cpu.rf_ram.memory[45][2] ),
    .A2(_02973_),
    .ZN(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07483_ (.A1(_02900_),
    .A2(_02969_),
    .B(_02974_),
    .ZN(_00116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07484_ (.A1(\u_cpu.rf_ram.memory[45][3] ),
    .A2(_02973_),
    .ZN(_02975_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07485_ (.A1(_02904_),
    .A2(_02969_),
    .B(_02975_),
    .ZN(_00117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07486_ (.A1(\u_cpu.rf_ram.memory[45][4] ),
    .A2(_02973_),
    .ZN(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07487_ (.A1(_02907_),
    .A2(_02969_),
    .B(_02976_),
    .ZN(_00118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07488_ (.A1(\u_cpu.rf_ram.memory[45][5] ),
    .A2(_02973_),
    .ZN(_02977_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07489_ (.A1(_02910_),
    .A2(_02970_),
    .B(_02977_),
    .ZN(_00119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07490_ (.A1(\u_cpu.rf_ram.memory[45][6] ),
    .A2(_02973_),
    .ZN(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07491_ (.A1(_02913_),
    .A2(_02970_),
    .B(_02978_),
    .ZN(_00120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07492_ (.A1(\u_cpu.rf_ram.memory[45][7] ),
    .A2(_02968_),
    .ZN(_02979_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07493_ (.A1(_02916_),
    .A2(_02970_),
    .B(_02979_),
    .ZN(_00121_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07494_ (.I(_02888_),
    .Z(_02980_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07495_ (.A1(_02829_),
    .A2(_02919_),
    .ZN(_02981_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07496_ (.I(_02981_),
    .Z(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07497_ (.A1(_02965_),
    .A2(_02982_),
    .ZN(_02983_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07498_ (.I(_02983_),
    .Z(_02984_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07499_ (.I(_02983_),
    .Z(_02985_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07500_ (.A1(\u_cpu.rf_ram.memory[44][0] ),
    .A2(_02985_),
    .ZN(_02986_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07501_ (.A1(_02980_),
    .A2(_02984_),
    .B(_02986_),
    .ZN(_00122_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07502_ (.I(_02896_),
    .Z(_02987_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07503_ (.A1(\u_cpu.rf_ram.memory[44][1] ),
    .A2(_02985_),
    .ZN(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07504_ (.A1(_02987_),
    .A2(_02984_),
    .B(_02988_),
    .ZN(_00123_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07505_ (.I(_02899_),
    .Z(_02989_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07506_ (.I(_02983_),
    .Z(_02990_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07507_ (.A1(\u_cpu.rf_ram.memory[44][2] ),
    .A2(_02990_),
    .ZN(_02991_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07508_ (.A1(_02989_),
    .A2(_02984_),
    .B(_02991_),
    .ZN(_00124_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07509_ (.I(_02903_),
    .Z(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07510_ (.A1(\u_cpu.rf_ram.memory[44][3] ),
    .A2(_02990_),
    .ZN(_02993_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07511_ (.A1(_02992_),
    .A2(_02984_),
    .B(_02993_),
    .ZN(_00125_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07512_ (.I(_02906_),
    .Z(_02994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07513_ (.A1(\u_cpu.rf_ram.memory[44][4] ),
    .A2(_02990_),
    .ZN(_02995_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07514_ (.A1(_02994_),
    .A2(_02984_),
    .B(_02995_),
    .ZN(_00126_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07515_ (.I(_02909_),
    .Z(_02996_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07516_ (.A1(\u_cpu.rf_ram.memory[44][5] ),
    .A2(_02990_),
    .ZN(_02997_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07517_ (.A1(_02996_),
    .A2(_02985_),
    .B(_02997_),
    .ZN(_00127_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07518_ (.I(_02912_),
    .Z(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07519_ (.A1(\u_cpu.rf_ram.memory[44][6] ),
    .A2(_02990_),
    .ZN(_02999_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07520_ (.A1(_02998_),
    .A2(_02985_),
    .B(_02999_),
    .ZN(_00128_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07521_ (.I(_02915_),
    .Z(_03000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07522_ (.A1(\u_cpu.rf_ram.memory[44][7] ),
    .A2(_02983_),
    .ZN(_03001_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07523_ (.A1(_03000_),
    .A2(_02985_),
    .B(_03001_),
    .ZN(_00129_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07524_ (.A1(_02716_),
    .A2(_02875_),
    .ZN(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07525_ (.A1(\u_cpu.cpu.immdec.imm11_7[2] ),
    .A2(\u_cpu.cpu.immdec.imm11_7[3] ),
    .A3(_02724_),
    .ZN(_03003_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07526_ (.A1(_02788_),
    .A2(_03003_),
    .ZN(_03004_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07527_ (.I(_03004_),
    .Z(_03005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07528_ (.A1(_03002_),
    .A2(_03005_),
    .ZN(_03006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07529_ (.I(_03006_),
    .Z(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07530_ (.I(_03006_),
    .Z(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07531_ (.A1(\u_cpu.rf_ram.memory[51][0] ),
    .A2(_03008_),
    .ZN(_03009_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07532_ (.A1(_02980_),
    .A2(_03007_),
    .B(_03009_),
    .ZN(_00130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07533_ (.A1(\u_cpu.rf_ram.memory[51][1] ),
    .A2(_03008_),
    .ZN(_03010_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07534_ (.A1(_02987_),
    .A2(_03007_),
    .B(_03010_),
    .ZN(_00131_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07535_ (.I(_03006_),
    .Z(_03011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07536_ (.A1(\u_cpu.rf_ram.memory[51][2] ),
    .A2(_03011_),
    .ZN(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07537_ (.A1(_02989_),
    .A2(_03007_),
    .B(_03012_),
    .ZN(_00132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07538_ (.A1(\u_cpu.rf_ram.memory[51][3] ),
    .A2(_03011_),
    .ZN(_03013_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07539_ (.A1(_02992_),
    .A2(_03007_),
    .B(_03013_),
    .ZN(_00133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07540_ (.A1(\u_cpu.rf_ram.memory[51][4] ),
    .A2(_03011_),
    .ZN(_03014_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07541_ (.A1(_02994_),
    .A2(_03007_),
    .B(_03014_),
    .ZN(_00134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07542_ (.A1(\u_cpu.rf_ram.memory[51][5] ),
    .A2(_03011_),
    .ZN(_03015_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07543_ (.A1(_02996_),
    .A2(_03008_),
    .B(_03015_),
    .ZN(_00135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07544_ (.A1(\u_cpu.rf_ram.memory[51][6] ),
    .A2(_03011_),
    .ZN(_03016_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07545_ (.A1(_02998_),
    .A2(_03008_),
    .B(_03016_),
    .ZN(_00136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07546_ (.A1(\u_cpu.rf_ram.memory[51][7] ),
    .A2(_03006_),
    .ZN(_03017_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07547_ (.A1(_03000_),
    .A2(_03008_),
    .B(_03017_),
    .ZN(_00137_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07548_ (.I(_02939_),
    .Z(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07549_ (.A1(_02782_),
    .A2(_02936_),
    .ZN(_03019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07550_ (.I(_03019_),
    .Z(_03020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07551_ (.A1(_03018_),
    .A2(_03020_),
    .ZN(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07552_ (.I(_03021_),
    .Z(_03022_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07553_ (.I(_03021_),
    .Z(_03023_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07554_ (.A1(\u_cpu.rf_ram.memory[41][0] ),
    .A2(_03023_),
    .ZN(_03024_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07555_ (.A1(_02980_),
    .A2(_03022_),
    .B(_03024_),
    .ZN(_00138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07556_ (.A1(\u_cpu.rf_ram.memory[41][1] ),
    .A2(_03023_),
    .ZN(_03025_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07557_ (.A1(_02987_),
    .A2(_03022_),
    .B(_03025_),
    .ZN(_00139_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07558_ (.I(_03021_),
    .Z(_03026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07559_ (.A1(\u_cpu.rf_ram.memory[41][2] ),
    .A2(_03026_),
    .ZN(_03027_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07560_ (.A1(_02989_),
    .A2(_03022_),
    .B(_03027_),
    .ZN(_00140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07561_ (.A1(\u_cpu.rf_ram.memory[41][3] ),
    .A2(_03026_),
    .ZN(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07562_ (.A1(_02992_),
    .A2(_03022_),
    .B(_03028_),
    .ZN(_00141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07563_ (.A1(\u_cpu.rf_ram.memory[41][4] ),
    .A2(_03026_),
    .ZN(_03029_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07564_ (.A1(_02994_),
    .A2(_03022_),
    .B(_03029_),
    .ZN(_00142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07565_ (.A1(\u_cpu.rf_ram.memory[41][5] ),
    .A2(_03026_),
    .ZN(_03030_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07566_ (.A1(_02996_),
    .A2(_03023_),
    .B(_03030_),
    .ZN(_00143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07567_ (.A1(\u_cpu.rf_ram.memory[41][6] ),
    .A2(_03026_),
    .ZN(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07568_ (.A1(_02998_),
    .A2(_03023_),
    .B(_03031_),
    .ZN(_00144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07569_ (.A1(\u_cpu.rf_ram.memory[41][7] ),
    .A2(_03021_),
    .ZN(_03032_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07570_ (.A1(_03000_),
    .A2(_03023_),
    .B(_03032_),
    .ZN(_00145_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07571_ (.A1(_02875_),
    .A2(_02936_),
    .ZN(_03033_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07572_ (.I(_03033_),
    .Z(_03034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07573_ (.A1(_03018_),
    .A2(_03034_),
    .ZN(_03035_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07574_ (.I(_03035_),
    .Z(_03036_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07575_ (.I(_03035_),
    .Z(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07576_ (.A1(\u_cpu.rf_ram.memory[43][0] ),
    .A2(_03037_),
    .ZN(_03038_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07577_ (.A1(_02980_),
    .A2(_03036_),
    .B(_03038_),
    .ZN(_00146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07578_ (.A1(\u_cpu.rf_ram.memory[43][1] ),
    .A2(_03037_),
    .ZN(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07579_ (.A1(_02987_),
    .A2(_03036_),
    .B(_03039_),
    .ZN(_00147_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07580_ (.I(_03035_),
    .Z(_03040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07581_ (.A1(\u_cpu.rf_ram.memory[43][2] ),
    .A2(_03040_),
    .ZN(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07582_ (.A1(_02989_),
    .A2(_03036_),
    .B(_03041_),
    .ZN(_00148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07583_ (.A1(\u_cpu.rf_ram.memory[43][3] ),
    .A2(_03040_),
    .ZN(_03042_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07584_ (.A1(_02992_),
    .A2(_03036_),
    .B(_03042_),
    .ZN(_00149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07585_ (.A1(\u_cpu.rf_ram.memory[43][4] ),
    .A2(_03040_),
    .ZN(_03043_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07586_ (.A1(_02994_),
    .A2(_03036_),
    .B(_03043_),
    .ZN(_00150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07587_ (.A1(\u_cpu.rf_ram.memory[43][5] ),
    .A2(_03040_),
    .ZN(_03044_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07588_ (.A1(_02996_),
    .A2(_03037_),
    .B(_03044_),
    .ZN(_00151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07589_ (.A1(\u_cpu.rf_ram.memory[43][6] ),
    .A2(_03040_),
    .ZN(_03045_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07590_ (.A1(_02998_),
    .A2(_03037_),
    .B(_03045_),
    .ZN(_00152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07591_ (.A1(\u_cpu.rf_ram.memory[43][7] ),
    .A2(_03035_),
    .ZN(_03046_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07592_ (.A1(_03000_),
    .A2(_03037_),
    .B(_03046_),
    .ZN(_00153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07593_ (.A1(_02891_),
    .A2(_03005_),
    .ZN(_03047_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07594_ (.I(_03047_),
    .Z(_03048_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07595_ (.I(_03047_),
    .Z(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07596_ (.A1(\u_cpu.rf_ram.memory[48][0] ),
    .A2(_03049_),
    .ZN(_03050_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07597_ (.A1(_02980_),
    .A2(_03048_),
    .B(_03050_),
    .ZN(_00154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07598_ (.A1(\u_cpu.rf_ram.memory[48][1] ),
    .A2(_03049_),
    .ZN(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07599_ (.A1(_02987_),
    .A2(_03048_),
    .B(_03051_),
    .ZN(_00155_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07600_ (.I(_03047_),
    .Z(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07601_ (.A1(\u_cpu.rf_ram.memory[48][2] ),
    .A2(_03052_),
    .ZN(_03053_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07602_ (.A1(_02989_),
    .A2(_03048_),
    .B(_03053_),
    .ZN(_00156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07603_ (.A1(\u_cpu.rf_ram.memory[48][3] ),
    .A2(_03052_),
    .ZN(_03054_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07604_ (.A1(_02992_),
    .A2(_03048_),
    .B(_03054_),
    .ZN(_00157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07605_ (.A1(\u_cpu.rf_ram.memory[48][4] ),
    .A2(_03052_),
    .ZN(_03055_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07606_ (.A1(_02994_),
    .A2(_03048_),
    .B(_03055_),
    .ZN(_00158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07607_ (.A1(\u_cpu.rf_ram.memory[48][5] ),
    .A2(_03052_),
    .ZN(_03056_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07608_ (.A1(_02996_),
    .A2(_03049_),
    .B(_03056_),
    .ZN(_00159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07609_ (.A1(\u_cpu.rf_ram.memory[48][6] ),
    .A2(_03052_),
    .ZN(_03057_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07610_ (.A1(_02998_),
    .A2(_03049_),
    .B(_03057_),
    .ZN(_00160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07611_ (.A1(\u_cpu.rf_ram.memory[48][7] ),
    .A2(_03047_),
    .ZN(_03058_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07612_ (.A1(_03000_),
    .A2(_03049_),
    .B(_03058_),
    .ZN(_00161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07613_ (.I(_02739_),
    .Z(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07614_ (.I(_03059_),
    .Z(_03060_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07615_ (.A1(_02875_),
    .A2(_02919_),
    .ZN(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07616_ (.I(_03061_),
    .Z(_03062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07617_ (.A1(_03018_),
    .A2(_03062_),
    .ZN(_03063_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07618_ (.I(_03063_),
    .Z(_03064_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07619_ (.I(_03063_),
    .Z(_03065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07620_ (.A1(\u_cpu.rf_ram.memory[47][0] ),
    .A2(_03065_),
    .ZN(_03066_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07621_ (.A1(_03060_),
    .A2(_03064_),
    .B(_03066_),
    .ZN(_00162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07622_ (.I(_02745_),
    .Z(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07623_ (.I(_03067_),
    .Z(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07624_ (.A1(\u_cpu.rf_ram.memory[47][1] ),
    .A2(_03065_),
    .ZN(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07625_ (.A1(_03068_),
    .A2(_03064_),
    .B(_03069_),
    .ZN(_00163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07626_ (.I(_02751_),
    .Z(_03070_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07627_ (.I(_03070_),
    .Z(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07628_ (.I(_03063_),
    .Z(_03072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07629_ (.A1(\u_cpu.rf_ram.memory[47][2] ),
    .A2(_03072_),
    .ZN(_03073_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07630_ (.A1(_03071_),
    .A2(_03064_),
    .B(_03073_),
    .ZN(_00164_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07631_ (.I(_02757_),
    .Z(_03074_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07632_ (.I(_03074_),
    .Z(_03075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07633_ (.A1(\u_cpu.rf_ram.memory[47][3] ),
    .A2(_03072_),
    .ZN(_03076_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07634_ (.A1(_03075_),
    .A2(_03064_),
    .B(_03076_),
    .ZN(_00165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07635_ (.I(_02762_),
    .Z(_03077_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07636_ (.I(_03077_),
    .Z(_03078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07637_ (.A1(\u_cpu.rf_ram.memory[47][4] ),
    .A2(_03072_),
    .ZN(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07638_ (.A1(_03078_),
    .A2(_03064_),
    .B(_03079_),
    .ZN(_00166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07639_ (.I(_02767_),
    .Z(_03080_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07640_ (.I(_03080_),
    .Z(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07641_ (.A1(\u_cpu.rf_ram.memory[47][5] ),
    .A2(_03072_),
    .ZN(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07642_ (.A1(_03081_),
    .A2(_03065_),
    .B(_03082_),
    .ZN(_00167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07643_ (.I(_02772_),
    .Z(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07644_ (.I(_03083_),
    .Z(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07645_ (.A1(\u_cpu.rf_ram.memory[47][6] ),
    .A2(_03072_),
    .ZN(_03085_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07646_ (.A1(_03084_),
    .A2(_03065_),
    .B(_03085_),
    .ZN(_00168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07647_ (.I(_02777_),
    .Z(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07648_ (.I(_03086_),
    .Z(_03087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07649_ (.A1(\u_cpu.rf_ram.memory[47][7] ),
    .A2(_03063_),
    .ZN(_03088_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07650_ (.A1(_03087_),
    .A2(_03065_),
    .B(_03088_),
    .ZN(_00169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07651_ (.A1(_02723_),
    .A2(_03005_),
    .ZN(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07652_ (.I(_03089_),
    .Z(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07653_ (.I(_03089_),
    .Z(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07654_ (.A1(\u_cpu.rf_ram.memory[50][0] ),
    .A2(_03091_),
    .ZN(_03092_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07655_ (.A1(_03060_),
    .A2(_03090_),
    .B(_03092_),
    .ZN(_00170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07656_ (.A1(\u_cpu.rf_ram.memory[50][1] ),
    .A2(_03091_),
    .ZN(_03093_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07657_ (.A1(_03068_),
    .A2(_03090_),
    .B(_03093_),
    .ZN(_00171_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07658_ (.I(_03089_),
    .Z(_03094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07659_ (.A1(\u_cpu.rf_ram.memory[50][2] ),
    .A2(_03094_),
    .ZN(_03095_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07660_ (.A1(_03071_),
    .A2(_03090_),
    .B(_03095_),
    .ZN(_00172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07661_ (.A1(\u_cpu.rf_ram.memory[50][3] ),
    .A2(_03094_),
    .ZN(_03096_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07662_ (.A1(_03075_),
    .A2(_03090_),
    .B(_03096_),
    .ZN(_00173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07663_ (.A1(\u_cpu.rf_ram.memory[50][4] ),
    .A2(_03094_),
    .ZN(_03097_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07664_ (.A1(_03078_),
    .A2(_03090_),
    .B(_03097_),
    .ZN(_00174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07665_ (.A1(\u_cpu.rf_ram.memory[50][5] ),
    .A2(_03094_),
    .ZN(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07666_ (.A1(_03081_),
    .A2(_03091_),
    .B(_03098_),
    .ZN(_00175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07667_ (.A1(\u_cpu.rf_ram.memory[50][6] ),
    .A2(_03094_),
    .ZN(_03099_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07668_ (.A1(_03084_),
    .A2(_03091_),
    .B(_03099_),
    .ZN(_00176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07669_ (.A1(\u_cpu.rf_ram.memory[50][7] ),
    .A2(_03089_),
    .ZN(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07670_ (.A1(_03087_),
    .A2(_03091_),
    .B(_03100_),
    .ZN(_00177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07671_ (.A1(_02831_),
    .A2(_02850_),
    .ZN(_03101_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07672_ (.I(_03101_),
    .Z(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07673_ (.I0(_02846_),
    .I1(\u_cpu.rf_ram.memory[4][0] ),
    .S(_03102_),
    .Z(_03103_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07674_ (.I(_03103_),
    .Z(_00178_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07675_ (.I0(_02855_),
    .I1(\u_cpu.rf_ram.memory[4][1] ),
    .S(_03102_),
    .Z(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07676_ (.I(_03104_),
    .Z(_00179_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07677_ (.I0(_02858_),
    .I1(\u_cpu.rf_ram.memory[4][2] ),
    .S(_03102_),
    .Z(_03105_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07678_ (.I(_03105_),
    .Z(_00180_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07679_ (.I0(_02861_),
    .I1(\u_cpu.rf_ram.memory[4][3] ),
    .S(_03102_),
    .Z(_03106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07680_ (.I(_03106_),
    .Z(_00181_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07681_ (.I0(_02864_),
    .I1(\u_cpu.rf_ram.memory[4][4] ),
    .S(_03102_),
    .Z(_03107_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07682_ (.I(_03107_),
    .Z(_00182_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07683_ (.I0(_02867_),
    .I1(\u_cpu.rf_ram.memory[4][5] ),
    .S(_03101_),
    .Z(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07684_ (.I(_03108_),
    .Z(_00183_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07685_ (.I0(_02870_),
    .I1(\u_cpu.rf_ram.memory[4][6] ),
    .S(_03101_),
    .Z(_03109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07686_ (.I(_03109_),
    .Z(_00184_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07687_ (.I0(_02873_),
    .I1(\u_cpu.rf_ram.memory[4][7] ),
    .S(_03101_),
    .Z(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07688_ (.I(_03110_),
    .Z(_00185_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07689_ (.I(net2),
    .Z(_03111_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07690_ (.I(_03111_),
    .Z(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07691_ (.I(_01437_),
    .ZN(_03113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07692_ (.I(_03113_),
    .Z(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07693_ (.I(_03114_),
    .Z(_03115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07694_ (.A1(net8),
    .A2(_01433_),
    .ZN(_03116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07695_ (.A1(_03115_),
    .A2(\u_arbiter.i_wb_cpu_ibus_adr[1] ),
    .B(_03116_),
    .ZN(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07696_ (.I(_03117_),
    .Z(_03118_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07697_ (.A1(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ),
    .A2(\u_cpu.cpu.state.stage_two_req ),
    .B(_03118_),
    .ZN(_03119_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07698_ (.A1(_03112_),
    .A2(_03119_),
    .ZN(_00186_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07699_ (.A1(_02569_),
    .A2(_02695_),
    .B(_02598_),
    .ZN(_03120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07700_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[6] ),
    .A2(_03120_),
    .ZN(_03121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07701_ (.A1(_01374_),
    .A2(_02556_),
    .ZN(_03122_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07702_ (.A1(_02694_),
    .A2(_02595_),
    .Z(_03123_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07703_ (.A1(_03122_),
    .A2(_03123_),
    .ZN(_03124_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07704_ (.I(\u_arbiter.i_wb_cpu_dbus_dat[0] ),
    .Z(_03125_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _07705_ (.A1(_03125_),
    .A2(net36),
    .A3(\u_arbiter.i_wb_cpu_dbus_dat[2] ),
    .A4(\u_arbiter.i_wb_cpu_dbus_dat[3] ),
    .Z(_03126_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07706_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[4] ),
    .A2(_03126_),
    .ZN(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07707_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .A2(_03127_),
    .Z(_03128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07708_ (.A1(_03124_),
    .A2(_03128_),
    .ZN(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07709_ (.A1(_03121_),
    .A2(_03129_),
    .ZN(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07710_ (.A1(_01409_),
    .A2(_02559_),
    .A3(_03130_),
    .ZN(_03131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07711_ (.A1(net8),
    .A2(_01450_),
    .ZN(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07712_ (.A1(_02605_),
    .A2(_03131_),
    .B(_03132_),
    .C(_02684_),
    .ZN(_03133_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _07713_ (.A1(_02597_),
    .A2(_01386_),
    .A3(_02674_),
    .A4(_03133_),
    .ZN(_03134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07714_ (.A1(_03119_),
    .A2(_03134_),
    .ZN(_03135_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07715_ (.A1(_02717_),
    .A2(_03135_),
    .ZN(_00187_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07716_ (.A1(\u_cpu.rf_ram_if.rcnt[2] ),
    .A2(\u_cpu.rf_ram_if.rcnt[1] ),
    .A3(_02717_),
    .Z(_03136_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07717_ (.A1(_02718_),
    .A2(_03135_),
    .A3(_03136_),
    .ZN(_00188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07718_ (.A1(_01820_),
    .A2(_03136_),
    .ZN(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07719_ (.A1(_01820_),
    .A2(_03136_),
    .Z(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _07720_ (.A1(_03119_),
    .A2(_03134_),
    .A3(_03137_),
    .A4(_03138_),
    .Z(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07721_ (.I(_03139_),
    .Z(_00189_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07722_ (.A1(_01821_),
    .A2(_03137_),
    .Z(_03140_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07723_ (.A1(_03135_),
    .A2(_03140_),
    .ZN(_00190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07724_ (.A1(_02790_),
    .A2(_02891_),
    .ZN(_03141_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07725_ (.I(_03141_),
    .Z(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07726_ (.I(_03141_),
    .Z(_03143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07727_ (.A1(\u_cpu.rf_ram.memory[16][0] ),
    .A2(_03143_),
    .ZN(_03144_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07728_ (.A1(_03060_),
    .A2(_03142_),
    .B(_03144_),
    .ZN(_00191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07729_ (.A1(\u_cpu.rf_ram.memory[16][1] ),
    .A2(_03143_),
    .ZN(_03145_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07730_ (.A1(_03068_),
    .A2(_03142_),
    .B(_03145_),
    .ZN(_00192_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07731_ (.I(_03141_),
    .Z(_03146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07732_ (.A1(\u_cpu.rf_ram.memory[16][2] ),
    .A2(_03146_),
    .ZN(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07733_ (.A1(_03071_),
    .A2(_03142_),
    .B(_03147_),
    .ZN(_00193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07734_ (.A1(\u_cpu.rf_ram.memory[16][3] ),
    .A2(_03146_),
    .ZN(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07735_ (.A1(_03075_),
    .A2(_03142_),
    .B(_03148_),
    .ZN(_00194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07736_ (.A1(\u_cpu.rf_ram.memory[16][4] ),
    .A2(_03146_),
    .ZN(_03149_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07737_ (.A1(_03078_),
    .A2(_03142_),
    .B(_03149_),
    .ZN(_00195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07738_ (.A1(\u_cpu.rf_ram.memory[16][5] ),
    .A2(_03146_),
    .ZN(_03150_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07739_ (.A1(_03081_),
    .A2(_03143_),
    .B(_03150_),
    .ZN(_00196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07740_ (.A1(\u_cpu.rf_ram.memory[16][6] ),
    .A2(_03146_),
    .ZN(_03151_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07741_ (.A1(_03084_),
    .A2(_03143_),
    .B(_03151_),
    .ZN(_00197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07742_ (.A1(\u_cpu.rf_ram.memory[16][7] ),
    .A2(_03141_),
    .ZN(_03152_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07743_ (.A1(_03087_),
    .A2(_03143_),
    .B(_03152_),
    .ZN(_00198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07744_ (.A1(_02790_),
    .A2(_02804_),
    .ZN(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07745_ (.I(_03153_),
    .Z(_03154_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07746_ (.I(_03153_),
    .Z(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07747_ (.A1(\u_cpu.rf_ram.memory[17][0] ),
    .A2(_03155_),
    .ZN(_03156_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07748_ (.A1(_03060_),
    .A2(_03154_),
    .B(_03156_),
    .ZN(_00199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07749_ (.A1(\u_cpu.rf_ram.memory[17][1] ),
    .A2(_03155_),
    .ZN(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07750_ (.A1(_03068_),
    .A2(_03154_),
    .B(_03157_),
    .ZN(_00200_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07751_ (.I(_03153_),
    .Z(_03158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07752_ (.A1(\u_cpu.rf_ram.memory[17][2] ),
    .A2(_03158_),
    .ZN(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07753_ (.A1(_03071_),
    .A2(_03154_),
    .B(_03159_),
    .ZN(_00201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07754_ (.A1(\u_cpu.rf_ram.memory[17][3] ),
    .A2(_03158_),
    .ZN(_03160_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07755_ (.A1(_03075_),
    .A2(_03154_),
    .B(_03160_),
    .ZN(_00202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07756_ (.A1(\u_cpu.rf_ram.memory[17][4] ),
    .A2(_03158_),
    .ZN(_03161_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07757_ (.A1(_03078_),
    .A2(_03154_),
    .B(_03161_),
    .ZN(_00203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07758_ (.A1(\u_cpu.rf_ram.memory[17][5] ),
    .A2(_03158_),
    .ZN(_03162_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07759_ (.A1(_03081_),
    .A2(_03155_),
    .B(_03162_),
    .ZN(_00204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07760_ (.A1(\u_cpu.rf_ram.memory[17][6] ),
    .A2(_03158_),
    .ZN(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07761_ (.A1(_03084_),
    .A2(_03155_),
    .B(_03163_),
    .ZN(_00205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07762_ (.A1(\u_cpu.rf_ram.memory[17][7] ),
    .A2(_03153_),
    .ZN(_03164_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07763_ (.A1(_03087_),
    .A2(_03155_),
    .B(_03164_),
    .ZN(_00206_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07764_ (.A1(_02829_),
    .A2(_02936_),
    .ZN(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07765_ (.I(_03165_),
    .Z(_03166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07766_ (.A1(_03018_),
    .A2(_03166_),
    .ZN(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07767_ (.I(_03167_),
    .Z(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07768_ (.I(_03167_),
    .Z(_03169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07769_ (.A1(\u_cpu.rf_ram.memory[40][0] ),
    .A2(_03169_),
    .ZN(_03170_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07770_ (.A1(_03060_),
    .A2(_03168_),
    .B(_03170_),
    .ZN(_00207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07771_ (.A1(\u_cpu.rf_ram.memory[40][1] ),
    .A2(_03169_),
    .ZN(_03171_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07772_ (.A1(_03068_),
    .A2(_03168_),
    .B(_03171_),
    .ZN(_00208_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07773_ (.I(_03167_),
    .Z(_03172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07774_ (.A1(\u_cpu.rf_ram.memory[40][2] ),
    .A2(_03172_),
    .ZN(_03173_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07775_ (.A1(_03071_),
    .A2(_03168_),
    .B(_03173_),
    .ZN(_00209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07776_ (.A1(\u_cpu.rf_ram.memory[40][3] ),
    .A2(_03172_),
    .ZN(_03174_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07777_ (.A1(_03075_),
    .A2(_03168_),
    .B(_03174_),
    .ZN(_00210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07778_ (.A1(\u_cpu.rf_ram.memory[40][4] ),
    .A2(_03172_),
    .ZN(_03175_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07779_ (.A1(_03078_),
    .A2(_03168_),
    .B(_03175_),
    .ZN(_00211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07780_ (.A1(\u_cpu.rf_ram.memory[40][5] ),
    .A2(_03172_),
    .ZN(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07781_ (.A1(_03081_),
    .A2(_03169_),
    .B(_03176_),
    .ZN(_00212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07782_ (.A1(\u_cpu.rf_ram.memory[40][6] ),
    .A2(_03172_),
    .ZN(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07783_ (.A1(_03084_),
    .A2(_03169_),
    .B(_03177_),
    .ZN(_00213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07784_ (.A1(\u_cpu.rf_ram.memory[40][7] ),
    .A2(_03167_),
    .ZN(_03178_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07785_ (.A1(_03087_),
    .A2(_03169_),
    .B(_03178_),
    .ZN(_00214_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07786_ (.I(_03059_),
    .Z(_03179_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07787_ (.A1(_02729_),
    .A2(_03003_),
    .ZN(_03180_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07788_ (.I(_03180_),
    .Z(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07789_ (.A1(_02877_),
    .A2(_03181_),
    .ZN(_03182_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07790_ (.I(_03182_),
    .Z(_03183_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07791_ (.I(_03182_),
    .Z(_03184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07792_ (.A1(\u_cpu.rf_ram.memory[119][0] ),
    .A2(_03184_),
    .ZN(_03185_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07793_ (.A1(_03179_),
    .A2(_03183_),
    .B(_03185_),
    .ZN(_00215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07794_ (.I(_03067_),
    .Z(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07795_ (.A1(\u_cpu.rf_ram.memory[119][1] ),
    .A2(_03184_),
    .ZN(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07796_ (.A1(_03186_),
    .A2(_03183_),
    .B(_03187_),
    .ZN(_00216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07797_ (.I(_03070_),
    .Z(_03188_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07798_ (.I(_03182_),
    .Z(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07799_ (.A1(\u_cpu.rf_ram.memory[119][2] ),
    .A2(_03189_),
    .ZN(_03190_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07800_ (.A1(_03188_),
    .A2(_03183_),
    .B(_03190_),
    .ZN(_00217_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07801_ (.I(_03074_),
    .Z(_03191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07802_ (.A1(\u_cpu.rf_ram.memory[119][3] ),
    .A2(_03189_),
    .ZN(_03192_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07803_ (.A1(_03191_),
    .A2(_03183_),
    .B(_03192_),
    .ZN(_00218_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07804_ (.I(_03077_),
    .Z(_03193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07805_ (.A1(\u_cpu.rf_ram.memory[119][4] ),
    .A2(_03189_),
    .ZN(_03194_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07806_ (.A1(_03193_),
    .A2(_03183_),
    .B(_03194_),
    .ZN(_00219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07807_ (.I(_03080_),
    .Z(_03195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07808_ (.A1(\u_cpu.rf_ram.memory[119][5] ),
    .A2(_03189_),
    .ZN(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07809_ (.A1(_03195_),
    .A2(_03184_),
    .B(_03196_),
    .ZN(_00220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07810_ (.I(_03083_),
    .Z(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07811_ (.A1(\u_cpu.rf_ram.memory[119][6] ),
    .A2(_03189_),
    .ZN(_03198_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07812_ (.A1(_03197_),
    .A2(_03184_),
    .B(_03198_),
    .ZN(_00221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07813_ (.I(_03086_),
    .Z(_03199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07814_ (.A1(\u_cpu.rf_ram.memory[119][7] ),
    .A2(_03182_),
    .ZN(_03200_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07815_ (.A1(_03199_),
    .A2(_03184_),
    .B(_03200_),
    .ZN(_00222_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07816_ (.A1(_02724_),
    .A2(_02727_),
    .ZN(_03201_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07817_ (.I(_03201_),
    .Z(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07818_ (.A1(_02804_),
    .A2(_03202_),
    .ZN(_03203_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07819_ (.I(_03203_),
    .Z(_03204_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07820_ (.I(_03203_),
    .Z(_03205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07821_ (.A1(\u_cpu.rf_ram.memory[129][0] ),
    .A2(_03205_),
    .ZN(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07822_ (.A1(_03179_),
    .A2(_03204_),
    .B(_03206_),
    .ZN(_00223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07823_ (.A1(\u_cpu.rf_ram.memory[129][1] ),
    .A2(_03205_),
    .ZN(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07824_ (.A1(_03186_),
    .A2(_03204_),
    .B(_03207_),
    .ZN(_00224_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07825_ (.I(_03203_),
    .Z(_03208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07826_ (.A1(\u_cpu.rf_ram.memory[129][2] ),
    .A2(_03208_),
    .ZN(_03209_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07827_ (.A1(_03188_),
    .A2(_03204_),
    .B(_03209_),
    .ZN(_00225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07828_ (.A1(\u_cpu.rf_ram.memory[129][3] ),
    .A2(_03208_),
    .ZN(_03210_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07829_ (.A1(_03191_),
    .A2(_03204_),
    .B(_03210_),
    .ZN(_00226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07830_ (.A1(\u_cpu.rf_ram.memory[129][4] ),
    .A2(_03208_),
    .ZN(_03211_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07831_ (.A1(_03193_),
    .A2(_03204_),
    .B(_03211_),
    .ZN(_00227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07832_ (.A1(\u_cpu.rf_ram.memory[129][5] ),
    .A2(_03208_),
    .ZN(_03212_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07833_ (.A1(_03195_),
    .A2(_03205_),
    .B(_03212_),
    .ZN(_00228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07834_ (.A1(\u_cpu.rf_ram.memory[129][6] ),
    .A2(_03208_),
    .ZN(_03213_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07835_ (.A1(_03197_),
    .A2(_03205_),
    .B(_03213_),
    .ZN(_00229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07836_ (.A1(\u_cpu.rf_ram.memory[129][7] ),
    .A2(_03203_),
    .ZN(_03214_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07837_ (.A1(_03199_),
    .A2(_03205_),
    .B(_03214_),
    .ZN(_00230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07838_ (.A1(_03033_),
    .A2(_03202_),
    .ZN(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07839_ (.I(_03215_),
    .Z(_03216_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07840_ (.I(_03215_),
    .Z(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07841_ (.A1(\u_cpu.rf_ram.memory[139][0] ),
    .A2(_03217_),
    .ZN(_03218_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07842_ (.A1(_03179_),
    .A2(_03216_),
    .B(_03218_),
    .ZN(_00231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07843_ (.A1(\u_cpu.rf_ram.memory[139][1] ),
    .A2(_03217_),
    .ZN(_03219_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07844_ (.A1(_03186_),
    .A2(_03216_),
    .B(_03219_),
    .ZN(_00232_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07845_ (.I(_03215_),
    .Z(_03220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07846_ (.A1(\u_cpu.rf_ram.memory[139][2] ),
    .A2(_03220_),
    .ZN(_03221_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07847_ (.A1(_03188_),
    .A2(_03216_),
    .B(_03221_),
    .ZN(_00233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07848_ (.A1(\u_cpu.rf_ram.memory[139][3] ),
    .A2(_03220_),
    .ZN(_03222_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07849_ (.A1(_03191_),
    .A2(_03216_),
    .B(_03222_),
    .ZN(_00234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07850_ (.A1(\u_cpu.rf_ram.memory[139][4] ),
    .A2(_03220_),
    .ZN(_03223_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07851_ (.A1(_03193_),
    .A2(_03216_),
    .B(_03223_),
    .ZN(_00235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07852_ (.A1(\u_cpu.rf_ram.memory[139][5] ),
    .A2(_03220_),
    .ZN(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07853_ (.A1(_03195_),
    .A2(_03217_),
    .B(_03224_),
    .ZN(_00236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07854_ (.A1(\u_cpu.rf_ram.memory[139][6] ),
    .A2(_03220_),
    .ZN(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07855_ (.A1(_03197_),
    .A2(_03217_),
    .B(_03225_),
    .ZN(_00237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07856_ (.A1(\u_cpu.rf_ram.memory[139][7] ),
    .A2(_03215_),
    .ZN(_03226_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07857_ (.A1(_03199_),
    .A2(_03217_),
    .B(_03226_),
    .ZN(_00238_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07858_ (.I(_02922_),
    .Z(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07859_ (.A1(_03227_),
    .A2(_02967_),
    .ZN(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07860_ (.I(_03228_),
    .Z(_03229_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07861_ (.I(_03228_),
    .Z(_03230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07862_ (.A1(\u_cpu.rf_ram.memory[77][0] ),
    .A2(_03230_),
    .ZN(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07863_ (.A1(_03179_),
    .A2(_03229_),
    .B(_03231_),
    .ZN(_00239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07864_ (.A1(\u_cpu.rf_ram.memory[77][1] ),
    .A2(_03230_),
    .ZN(_03232_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07865_ (.A1(_03186_),
    .A2(_03229_),
    .B(_03232_),
    .ZN(_00240_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07866_ (.I(_03228_),
    .Z(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07867_ (.A1(\u_cpu.rf_ram.memory[77][2] ),
    .A2(_03233_),
    .ZN(_03234_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07868_ (.A1(_03188_),
    .A2(_03229_),
    .B(_03234_),
    .ZN(_00241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07869_ (.A1(\u_cpu.rf_ram.memory[77][3] ),
    .A2(_03233_),
    .ZN(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07870_ (.A1(_03191_),
    .A2(_03229_),
    .B(_03235_),
    .ZN(_00242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07871_ (.A1(\u_cpu.rf_ram.memory[77][4] ),
    .A2(_03233_),
    .ZN(_03236_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07872_ (.A1(_03193_),
    .A2(_03229_),
    .B(_03236_),
    .ZN(_00243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07873_ (.A1(\u_cpu.rf_ram.memory[77][5] ),
    .A2(_03233_),
    .ZN(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07874_ (.A1(_03195_),
    .A2(_03230_),
    .B(_03237_),
    .ZN(_00244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07875_ (.A1(\u_cpu.rf_ram.memory[77][6] ),
    .A2(_03233_),
    .ZN(_03238_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07876_ (.A1(_03197_),
    .A2(_03230_),
    .B(_03238_),
    .ZN(_00245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07877_ (.A1(\u_cpu.rf_ram.memory[77][7] ),
    .A2(_03228_),
    .ZN(_03239_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07878_ (.A1(_03199_),
    .A2(_03230_),
    .B(_03239_),
    .ZN(_00246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07879_ (.A1(_03227_),
    .A2(_02938_),
    .ZN(_03240_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07880_ (.I(_03240_),
    .Z(_03241_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07881_ (.I(_03240_),
    .Z(_03242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07882_ (.A1(\u_cpu.rf_ram.memory[74][0] ),
    .A2(_03242_),
    .ZN(_03243_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07883_ (.A1(_03179_),
    .A2(_03241_),
    .B(_03243_),
    .ZN(_00247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07884_ (.A1(\u_cpu.rf_ram.memory[74][1] ),
    .A2(_03242_),
    .ZN(_03244_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07885_ (.A1(_03186_),
    .A2(_03241_),
    .B(_03244_),
    .ZN(_00248_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07886_ (.I(_03240_),
    .Z(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07887_ (.A1(\u_cpu.rf_ram.memory[74][2] ),
    .A2(_03245_),
    .ZN(_03246_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07888_ (.A1(_03188_),
    .A2(_03241_),
    .B(_03246_),
    .ZN(_00249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07889_ (.A1(\u_cpu.rf_ram.memory[74][3] ),
    .A2(_03245_),
    .ZN(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07890_ (.A1(_03191_),
    .A2(_03241_),
    .B(_03247_),
    .ZN(_00250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07891_ (.A1(\u_cpu.rf_ram.memory[74][4] ),
    .A2(_03245_),
    .ZN(_03248_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07892_ (.A1(_03193_),
    .A2(_03241_),
    .B(_03248_),
    .ZN(_00251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07893_ (.A1(\u_cpu.rf_ram.memory[74][5] ),
    .A2(_03245_),
    .ZN(_03249_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07894_ (.A1(_03195_),
    .A2(_03242_),
    .B(_03249_),
    .ZN(_00252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07895_ (.A1(\u_cpu.rf_ram.memory[74][6] ),
    .A2(_03245_),
    .ZN(_03250_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07896_ (.A1(_03197_),
    .A2(_03242_),
    .B(_03250_),
    .ZN(_00253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07897_ (.A1(\u_cpu.rf_ram.memory[74][7] ),
    .A2(_03240_),
    .ZN(_03251_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07898_ (.A1(_03199_),
    .A2(_03242_),
    .B(_03251_),
    .ZN(_00254_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07899_ (.I(_03059_),
    .Z(_03252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07900_ (.A1(_03227_),
    .A2(_02982_),
    .ZN(_03253_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07901_ (.I(_03253_),
    .Z(_03254_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07902_ (.I(_03253_),
    .Z(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07903_ (.A1(\u_cpu.rf_ram.memory[76][0] ),
    .A2(_03255_),
    .ZN(_03256_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07904_ (.A1(_03252_),
    .A2(_03254_),
    .B(_03256_),
    .ZN(_00255_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07905_ (.I(_03067_),
    .Z(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07906_ (.A1(\u_cpu.rf_ram.memory[76][1] ),
    .A2(_03255_),
    .ZN(_03258_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07907_ (.A1(_03257_),
    .A2(_03254_),
    .B(_03258_),
    .ZN(_00256_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07908_ (.I(_03070_),
    .Z(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07909_ (.I(_03253_),
    .Z(_03260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07910_ (.A1(\u_cpu.rf_ram.memory[76][2] ),
    .A2(_03260_),
    .ZN(_03261_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07911_ (.A1(_03259_),
    .A2(_03254_),
    .B(_03261_),
    .ZN(_00257_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07912_ (.I(_03074_),
    .Z(_03262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07913_ (.A1(\u_cpu.rf_ram.memory[76][3] ),
    .A2(_03260_),
    .ZN(_03263_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07914_ (.A1(_03262_),
    .A2(_03254_),
    .B(_03263_),
    .ZN(_00258_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07915_ (.I(_03077_),
    .Z(_03264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07916_ (.A1(\u_cpu.rf_ram.memory[76][4] ),
    .A2(_03260_),
    .ZN(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07917_ (.A1(_03264_),
    .A2(_03254_),
    .B(_03265_),
    .ZN(_00259_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07918_ (.I(_03080_),
    .Z(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07919_ (.A1(\u_cpu.rf_ram.memory[76][5] ),
    .A2(_03260_),
    .ZN(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07920_ (.A1(_03266_),
    .A2(_03255_),
    .B(_03267_),
    .ZN(_00260_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07921_ (.I(_03083_),
    .Z(_03268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07922_ (.A1(\u_cpu.rf_ram.memory[76][6] ),
    .A2(_03260_),
    .ZN(_03269_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07923_ (.A1(_03268_),
    .A2(_03255_),
    .B(_03269_),
    .ZN(_00261_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07924_ (.I(_03086_),
    .Z(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07925_ (.A1(\u_cpu.rf_ram.memory[76][7] ),
    .A2(_03253_),
    .ZN(_03271_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07926_ (.A1(_03270_),
    .A2(_03255_),
    .B(_03271_),
    .ZN(_00262_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07927_ (.I(_02922_),
    .Z(_03272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07928_ (.A1(_03272_),
    .A2(_03034_),
    .ZN(_03273_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07929_ (.I(_03273_),
    .Z(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07930_ (.I(_03273_),
    .Z(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07931_ (.A1(\u_cpu.rf_ram.memory[75][0] ),
    .A2(_03275_),
    .ZN(_03276_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07932_ (.A1(_03252_),
    .A2(_03274_),
    .B(_03276_),
    .ZN(_00263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07933_ (.A1(\u_cpu.rf_ram.memory[75][1] ),
    .A2(_03275_),
    .ZN(_03277_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07934_ (.A1(_03257_),
    .A2(_03274_),
    .B(_03277_),
    .ZN(_00264_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07935_ (.I(_03273_),
    .Z(_03278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07936_ (.A1(\u_cpu.rf_ram.memory[75][2] ),
    .A2(_03278_),
    .ZN(_03279_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07937_ (.A1(_03259_),
    .A2(_03274_),
    .B(_03279_),
    .ZN(_00265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07938_ (.A1(\u_cpu.rf_ram.memory[75][3] ),
    .A2(_03278_),
    .ZN(_03280_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07939_ (.A1(_03262_),
    .A2(_03274_),
    .B(_03280_),
    .ZN(_00266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07940_ (.A1(\u_cpu.rf_ram.memory[75][4] ),
    .A2(_03278_),
    .ZN(_03281_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07941_ (.A1(_03264_),
    .A2(_03274_),
    .B(_03281_),
    .ZN(_00267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07942_ (.A1(\u_cpu.rf_ram.memory[75][5] ),
    .A2(_03278_),
    .ZN(_03282_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07943_ (.A1(_03266_),
    .A2(_03275_),
    .B(_03282_),
    .ZN(_00268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07944_ (.A1(\u_cpu.rf_ram.memory[75][6] ),
    .A2(_03278_),
    .ZN(_03283_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07945_ (.A1(_03268_),
    .A2(_03275_),
    .B(_03283_),
    .ZN(_00269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07946_ (.A1(\u_cpu.rf_ram.memory[75][7] ),
    .A2(_03273_),
    .ZN(_03284_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07947_ (.A1(_03270_),
    .A2(_03275_),
    .B(_03284_),
    .ZN(_00270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07948_ (.I(_02849_),
    .Z(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07949_ (.A1(_02721_),
    .A2(_02784_),
    .ZN(_03286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07950_ (.I(_03286_),
    .Z(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07951_ (.A1(_03285_),
    .A2(_03287_),
    .ZN(_03288_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07952_ (.I(_03288_),
    .Z(_03289_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07953_ (.I0(_02846_),
    .I1(\u_cpu.rf_ram.memory[6][0] ),
    .S(_03289_),
    .Z(_03290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07954_ (.I(_03290_),
    .Z(_00271_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07955_ (.I0(_02855_),
    .I1(\u_cpu.rf_ram.memory[6][1] ),
    .S(_03289_),
    .Z(_03291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07956_ (.I(_03291_),
    .Z(_00272_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07957_ (.I0(_02858_),
    .I1(\u_cpu.rf_ram.memory[6][2] ),
    .S(_03289_),
    .Z(_03292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07958_ (.I(_03292_),
    .Z(_00273_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07959_ (.I0(_02861_),
    .I1(\u_cpu.rf_ram.memory[6][3] ),
    .S(_03289_),
    .Z(_03293_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07960_ (.I(_03293_),
    .Z(_00274_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07961_ (.I0(_02864_),
    .I1(\u_cpu.rf_ram.memory[6][4] ),
    .S(_03289_),
    .Z(_03294_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07962_ (.I(_03294_),
    .Z(_00275_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07963_ (.I0(_02867_),
    .I1(\u_cpu.rf_ram.memory[6][5] ),
    .S(_03288_),
    .Z(_03295_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07964_ (.I(_03295_),
    .Z(_00276_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07965_ (.I0(_02870_),
    .I1(\u_cpu.rf_ram.memory[6][6] ),
    .S(_03288_),
    .Z(_03296_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07966_ (.I(_03296_),
    .Z(_00277_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07967_ (.I0(_02873_),
    .I1(\u_cpu.rf_ram.memory[6][7] ),
    .S(_03288_),
    .Z(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07968_ (.I(_03297_),
    .Z(_00278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07969_ (.A1(_02831_),
    .A2(_02923_),
    .ZN(_03298_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07970_ (.I(_03298_),
    .Z(_03299_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07971_ (.I(_03298_),
    .Z(_03300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07972_ (.A1(\u_cpu.rf_ram.memory[68][0] ),
    .A2(_03300_),
    .ZN(_03301_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07973_ (.A1(_03252_),
    .A2(_03299_),
    .B(_03301_),
    .ZN(_00279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07974_ (.A1(\u_cpu.rf_ram.memory[68][1] ),
    .A2(_03300_),
    .ZN(_03302_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07975_ (.A1(_03257_),
    .A2(_03299_),
    .B(_03302_),
    .ZN(_00280_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07976_ (.I(_03298_),
    .Z(_03303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07977_ (.A1(\u_cpu.rf_ram.memory[68][2] ),
    .A2(_03303_),
    .ZN(_03304_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07978_ (.A1(_03259_),
    .A2(_03299_),
    .B(_03304_),
    .ZN(_00281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07979_ (.A1(\u_cpu.rf_ram.memory[68][3] ),
    .A2(_03303_),
    .ZN(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07980_ (.A1(_03262_),
    .A2(_03299_),
    .B(_03305_),
    .ZN(_00282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07981_ (.A1(\u_cpu.rf_ram.memory[68][4] ),
    .A2(_03303_),
    .ZN(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07982_ (.A1(_03264_),
    .A2(_03299_),
    .B(_03306_),
    .ZN(_00283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07983_ (.A1(\u_cpu.rf_ram.memory[68][5] ),
    .A2(_03303_),
    .ZN(_03307_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07984_ (.A1(_03266_),
    .A2(_03300_),
    .B(_03307_),
    .ZN(_00284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07985_ (.A1(\u_cpu.rf_ram.memory[68][6] ),
    .A2(_03303_),
    .ZN(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07986_ (.A1(_03268_),
    .A2(_03300_),
    .B(_03308_),
    .ZN(_00285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07987_ (.A1(\u_cpu.rf_ram.memory[68][7] ),
    .A2(_03298_),
    .ZN(_03309_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07988_ (.A1(_03270_),
    .A2(_03300_),
    .B(_03309_),
    .ZN(_00286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07989_ (.I(_03002_),
    .Z(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07990_ (.A1(_03272_),
    .A2(_03310_),
    .ZN(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07991_ (.I(_03311_),
    .Z(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07992_ (.I(_03311_),
    .Z(_03313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07993_ (.A1(\u_cpu.rf_ram.memory[67][0] ),
    .A2(_03313_),
    .ZN(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07994_ (.A1(_03252_),
    .A2(_03312_),
    .B(_03314_),
    .ZN(_00287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07995_ (.A1(\u_cpu.rf_ram.memory[67][1] ),
    .A2(_03313_),
    .ZN(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07996_ (.A1(_03257_),
    .A2(_03312_),
    .B(_03315_),
    .ZN(_00288_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07997_ (.I(_03311_),
    .Z(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07998_ (.A1(\u_cpu.rf_ram.memory[67][2] ),
    .A2(_03316_),
    .ZN(_03317_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07999_ (.A1(_03259_),
    .A2(_03312_),
    .B(_03317_),
    .ZN(_00289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08000_ (.A1(\u_cpu.rf_ram.memory[67][3] ),
    .A2(_03316_),
    .ZN(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08001_ (.A1(_03262_),
    .A2(_03312_),
    .B(_03318_),
    .ZN(_00290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08002_ (.A1(\u_cpu.rf_ram.memory[67][4] ),
    .A2(_03316_),
    .ZN(_03319_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08003_ (.A1(_03264_),
    .A2(_03312_),
    .B(_03319_),
    .ZN(_00291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08004_ (.A1(\u_cpu.rf_ram.memory[67][5] ),
    .A2(_03316_),
    .ZN(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08005_ (.A1(_03266_),
    .A2(_03313_),
    .B(_03320_),
    .ZN(_00292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08006_ (.A1(\u_cpu.rf_ram.memory[67][6] ),
    .A2(_03316_),
    .ZN(_03321_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08007_ (.A1(_03268_),
    .A2(_03313_),
    .B(_03321_),
    .ZN(_00293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08008_ (.A1(\u_cpu.rf_ram.memory[67][7] ),
    .A2(_03311_),
    .ZN(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08009_ (.A1(_03270_),
    .A2(_03313_),
    .B(_03322_),
    .ZN(_00294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08010_ (.A1(_02723_),
    .A2(_02923_),
    .ZN(_03323_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08011_ (.I(_03323_),
    .Z(_03324_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08012_ (.I(_03323_),
    .Z(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08013_ (.A1(\u_cpu.rf_ram.memory[66][0] ),
    .A2(_03325_),
    .ZN(_03326_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08014_ (.A1(_03252_),
    .A2(_03324_),
    .B(_03326_),
    .ZN(_00295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08015_ (.A1(\u_cpu.rf_ram.memory[66][1] ),
    .A2(_03325_),
    .ZN(_03327_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08016_ (.A1(_03257_),
    .A2(_03324_),
    .B(_03327_),
    .ZN(_00296_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08017_ (.I(_03323_),
    .Z(_03328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08018_ (.A1(\u_cpu.rf_ram.memory[66][2] ),
    .A2(_03328_),
    .ZN(_03329_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08019_ (.A1(_03259_),
    .A2(_03324_),
    .B(_03329_),
    .ZN(_00297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08020_ (.A1(\u_cpu.rf_ram.memory[66][3] ),
    .A2(_03328_),
    .ZN(_03330_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08021_ (.A1(_03262_),
    .A2(_03324_),
    .B(_03330_),
    .ZN(_00298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08022_ (.A1(\u_cpu.rf_ram.memory[66][4] ),
    .A2(_03328_),
    .ZN(_03331_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08023_ (.A1(_03264_),
    .A2(_03324_),
    .B(_03331_),
    .ZN(_00299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08024_ (.A1(\u_cpu.rf_ram.memory[66][5] ),
    .A2(_03328_),
    .ZN(_03332_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08025_ (.A1(_03266_),
    .A2(_03325_),
    .B(_03332_),
    .ZN(_00300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08026_ (.A1(\u_cpu.rf_ram.memory[66][6] ),
    .A2(_03328_),
    .ZN(_03333_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08027_ (.A1(_03268_),
    .A2(_03325_),
    .B(_03333_),
    .ZN(_00301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08028_ (.A1(\u_cpu.rf_ram.memory[66][7] ),
    .A2(_03323_),
    .ZN(_03334_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08029_ (.A1(_03270_),
    .A2(_03325_),
    .B(_03334_),
    .ZN(_00302_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08030_ (.I(_03059_),
    .Z(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08031_ (.A1(_02804_),
    .A2(_02923_),
    .ZN(_03336_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08032_ (.I(_03336_),
    .Z(_03337_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08033_ (.I(_03336_),
    .Z(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08034_ (.A1(\u_cpu.rf_ram.memory[65][0] ),
    .A2(_03338_),
    .ZN(_03339_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08035_ (.A1(_03335_),
    .A2(_03337_),
    .B(_03339_),
    .ZN(_00303_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08036_ (.I(_03067_),
    .Z(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08037_ (.A1(\u_cpu.rf_ram.memory[65][1] ),
    .A2(_03338_),
    .ZN(_03341_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08038_ (.A1(_03340_),
    .A2(_03337_),
    .B(_03341_),
    .ZN(_00304_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08039_ (.I(_03070_),
    .Z(_03342_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08040_ (.I(_03336_),
    .Z(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08041_ (.A1(\u_cpu.rf_ram.memory[65][2] ),
    .A2(_03343_),
    .ZN(_03344_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08042_ (.A1(_03342_),
    .A2(_03337_),
    .B(_03344_),
    .ZN(_00305_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08043_ (.I(_03074_),
    .Z(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08044_ (.A1(\u_cpu.rf_ram.memory[65][3] ),
    .A2(_03343_),
    .ZN(_03346_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08045_ (.A1(_03345_),
    .A2(_03337_),
    .B(_03346_),
    .ZN(_00306_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08046_ (.I(_03077_),
    .Z(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08047_ (.A1(\u_cpu.rf_ram.memory[65][4] ),
    .A2(_03343_),
    .ZN(_03348_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08048_ (.A1(_03347_),
    .A2(_03337_),
    .B(_03348_),
    .ZN(_00307_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08049_ (.I(_03080_),
    .Z(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08050_ (.A1(\u_cpu.rf_ram.memory[65][5] ),
    .A2(_03343_),
    .ZN(_03350_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08051_ (.A1(_03349_),
    .A2(_03338_),
    .B(_03350_),
    .ZN(_00308_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08052_ (.I(_03083_),
    .Z(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08053_ (.A1(\u_cpu.rf_ram.memory[65][6] ),
    .A2(_03343_),
    .ZN(_03352_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08054_ (.A1(_03351_),
    .A2(_03338_),
    .B(_03352_),
    .ZN(_00309_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08055_ (.I(_03086_),
    .Z(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08056_ (.A1(\u_cpu.rf_ram.memory[65][7] ),
    .A2(_03336_),
    .ZN(_03354_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08057_ (.A1(_03353_),
    .A2(_03338_),
    .B(_03354_),
    .ZN(_00310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08058_ (.A1(_02891_),
    .A2(_02923_),
    .ZN(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08059_ (.I(_03355_),
    .Z(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08060_ (.I(_03355_),
    .Z(_03357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08061_ (.A1(\u_cpu.rf_ram.memory[64][0] ),
    .A2(_03357_),
    .ZN(_03358_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08062_ (.A1(_03335_),
    .A2(_03356_),
    .B(_03358_),
    .ZN(_00311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08063_ (.A1(\u_cpu.rf_ram.memory[64][1] ),
    .A2(_03357_),
    .ZN(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08064_ (.A1(_03340_),
    .A2(_03356_),
    .B(_03359_),
    .ZN(_00312_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08065_ (.I(_03355_),
    .Z(_03360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08066_ (.A1(\u_cpu.rf_ram.memory[64][2] ),
    .A2(_03360_),
    .ZN(_03361_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08067_ (.A1(_03342_),
    .A2(_03356_),
    .B(_03361_),
    .ZN(_00313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08068_ (.A1(\u_cpu.rf_ram.memory[64][3] ),
    .A2(_03360_),
    .ZN(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08069_ (.A1(_03345_),
    .A2(_03356_),
    .B(_03362_),
    .ZN(_00314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08070_ (.A1(\u_cpu.rf_ram.memory[64][4] ),
    .A2(_03360_),
    .ZN(_03363_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08071_ (.A1(_03347_),
    .A2(_03356_),
    .B(_03363_),
    .ZN(_00315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08072_ (.A1(\u_cpu.rf_ram.memory[64][5] ),
    .A2(_03360_),
    .ZN(_03364_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08073_ (.A1(_03349_),
    .A2(_03357_),
    .B(_03364_),
    .ZN(_00316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08074_ (.A1(\u_cpu.rf_ram.memory[64][6] ),
    .A2(_03360_),
    .ZN(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08075_ (.A1(_03351_),
    .A2(_03357_),
    .B(_03365_),
    .ZN(_00317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08076_ (.A1(\u_cpu.rf_ram.memory[64][7] ),
    .A2(_03355_),
    .ZN(_03366_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08077_ (.A1(_03353_),
    .A2(_03357_),
    .B(_03366_),
    .ZN(_00318_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08078_ (.I(_02789_),
    .Z(_03367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08079_ (.A1(_03367_),
    .A2(_02967_),
    .ZN(_03368_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08080_ (.I(_03368_),
    .Z(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08081_ (.I(_03368_),
    .Z(_03370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08082_ (.A1(\u_cpu.rf_ram.memory[29][0] ),
    .A2(_03370_),
    .ZN(_03371_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08083_ (.A1(_03335_),
    .A2(_03369_),
    .B(_03371_),
    .ZN(_00319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08084_ (.A1(\u_cpu.rf_ram.memory[29][1] ),
    .A2(_03370_),
    .ZN(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08085_ (.A1(_03340_),
    .A2(_03369_),
    .B(_03372_),
    .ZN(_00320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08086_ (.I(_03368_),
    .Z(_03373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08087_ (.A1(\u_cpu.rf_ram.memory[29][2] ),
    .A2(_03373_),
    .ZN(_03374_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08088_ (.A1(_03342_),
    .A2(_03369_),
    .B(_03374_),
    .ZN(_00321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08089_ (.A1(\u_cpu.rf_ram.memory[29][3] ),
    .A2(_03373_),
    .ZN(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08090_ (.A1(_03345_),
    .A2(_03369_),
    .B(_03375_),
    .ZN(_00322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08091_ (.A1(\u_cpu.rf_ram.memory[29][4] ),
    .A2(_03373_),
    .ZN(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08092_ (.A1(_03347_),
    .A2(_03369_),
    .B(_03376_),
    .ZN(_00323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08093_ (.A1(\u_cpu.rf_ram.memory[29][5] ),
    .A2(_03373_),
    .ZN(_03377_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08094_ (.A1(_03349_),
    .A2(_03370_),
    .B(_03377_),
    .ZN(_00324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08095_ (.A1(\u_cpu.rf_ram.memory[29][6] ),
    .A2(_03373_),
    .ZN(_03378_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08096_ (.A1(_03351_),
    .A2(_03370_),
    .B(_03378_),
    .ZN(_00325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08097_ (.A1(\u_cpu.rf_ram.memory[29][7] ),
    .A2(_03368_),
    .ZN(_03379_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08098_ (.A1(_03353_),
    .A2(_03370_),
    .B(_03379_),
    .ZN(_00326_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08099_ (.I(_03004_),
    .Z(_03380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08100_ (.A1(_03380_),
    .A2(_03062_),
    .ZN(_03381_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08101_ (.I(_03381_),
    .Z(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08102_ (.I(_03381_),
    .Z(_03383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08103_ (.A1(\u_cpu.rf_ram.memory[63][0] ),
    .A2(_03383_),
    .ZN(_03384_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08104_ (.A1(_03335_),
    .A2(_03382_),
    .B(_03384_),
    .ZN(_00327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08105_ (.A1(\u_cpu.rf_ram.memory[63][1] ),
    .A2(_03383_),
    .ZN(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08106_ (.A1(_03340_),
    .A2(_03382_),
    .B(_03385_),
    .ZN(_00328_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08107_ (.I(_03381_),
    .Z(_03386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08108_ (.A1(\u_cpu.rf_ram.memory[63][2] ),
    .A2(_03386_),
    .ZN(_03387_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08109_ (.A1(_03342_),
    .A2(_03382_),
    .B(_03387_),
    .ZN(_00329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08110_ (.A1(\u_cpu.rf_ram.memory[63][3] ),
    .A2(_03386_),
    .ZN(_03388_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08111_ (.A1(_03345_),
    .A2(_03382_),
    .B(_03388_),
    .ZN(_00330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08112_ (.A1(\u_cpu.rf_ram.memory[63][4] ),
    .A2(_03386_),
    .ZN(_03389_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08113_ (.A1(_03347_),
    .A2(_03382_),
    .B(_03389_),
    .ZN(_00331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08114_ (.A1(\u_cpu.rf_ram.memory[63][5] ),
    .A2(_03386_),
    .ZN(_03390_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08115_ (.A1(_03349_),
    .A2(_03383_),
    .B(_03390_),
    .ZN(_00332_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08116_ (.A1(\u_cpu.rf_ram.memory[63][6] ),
    .A2(_03386_),
    .ZN(_03391_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08117_ (.A1(_03351_),
    .A2(_03383_),
    .B(_03391_),
    .ZN(_00333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08118_ (.A1(\u_cpu.rf_ram.memory[63][7] ),
    .A2(_03381_),
    .ZN(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08119_ (.A1(_03353_),
    .A2(_03383_),
    .B(_03392_),
    .ZN(_00334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08120_ (.A1(_02920_),
    .A2(_03005_),
    .ZN(_03393_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08121_ (.I(_03393_),
    .Z(_03394_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08122_ (.I(_03393_),
    .Z(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08123_ (.A1(\u_cpu.rf_ram.memory[62][0] ),
    .A2(_03395_),
    .ZN(_03396_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08124_ (.A1(_03335_),
    .A2(_03394_),
    .B(_03396_),
    .ZN(_00335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08125_ (.A1(\u_cpu.rf_ram.memory[62][1] ),
    .A2(_03395_),
    .ZN(_03397_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08126_ (.A1(_03340_),
    .A2(_03394_),
    .B(_03397_),
    .ZN(_00336_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08127_ (.I(_03393_),
    .Z(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08128_ (.A1(\u_cpu.rf_ram.memory[62][2] ),
    .A2(_03398_),
    .ZN(_03399_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08129_ (.A1(_03342_),
    .A2(_03394_),
    .B(_03399_),
    .ZN(_00337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08130_ (.A1(\u_cpu.rf_ram.memory[62][3] ),
    .A2(_03398_),
    .ZN(_03400_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08131_ (.A1(_03345_),
    .A2(_03394_),
    .B(_03400_),
    .ZN(_00338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08132_ (.A1(\u_cpu.rf_ram.memory[62][4] ),
    .A2(_03398_),
    .ZN(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08133_ (.A1(_03347_),
    .A2(_03394_),
    .B(_03401_),
    .ZN(_00339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08134_ (.A1(\u_cpu.rf_ram.memory[62][5] ),
    .A2(_03398_),
    .ZN(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08135_ (.A1(_03349_),
    .A2(_03395_),
    .B(_03402_),
    .ZN(_00340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08136_ (.A1(\u_cpu.rf_ram.memory[62][6] ),
    .A2(_03398_),
    .ZN(_03403_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08137_ (.A1(_03351_),
    .A2(_03395_),
    .B(_03403_),
    .ZN(_00341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08138_ (.A1(\u_cpu.rf_ram.memory[62][7] ),
    .A2(_03393_),
    .ZN(_03404_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08139_ (.A1(_03353_),
    .A2(_03395_),
    .B(_03404_),
    .ZN(_00342_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08140_ (.I(_03059_),
    .Z(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08141_ (.A1(_02966_),
    .A2(_03005_),
    .ZN(_03406_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08142_ (.I(_03406_),
    .Z(_03407_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08143_ (.I(_03406_),
    .Z(_03408_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08144_ (.A1(\u_cpu.rf_ram.memory[61][0] ),
    .A2(_03408_),
    .ZN(_03409_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08145_ (.A1(_03405_),
    .A2(_03407_),
    .B(_03409_),
    .ZN(_00343_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08146_ (.I(_03067_),
    .Z(_03410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08147_ (.A1(\u_cpu.rf_ram.memory[61][1] ),
    .A2(_03408_),
    .ZN(_03411_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08148_ (.A1(_03410_),
    .A2(_03407_),
    .B(_03411_),
    .ZN(_00344_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08149_ (.I(_03070_),
    .Z(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08150_ (.I(_03406_),
    .Z(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08151_ (.A1(\u_cpu.rf_ram.memory[61][2] ),
    .A2(_03413_),
    .ZN(_03414_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08152_ (.A1(_03412_),
    .A2(_03407_),
    .B(_03414_),
    .ZN(_00345_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08153_ (.I(_03074_),
    .Z(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08154_ (.A1(\u_cpu.rf_ram.memory[61][3] ),
    .A2(_03413_),
    .ZN(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08155_ (.A1(_03415_),
    .A2(_03407_),
    .B(_03416_),
    .ZN(_00346_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08156_ (.I(_03077_),
    .Z(_03417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08157_ (.A1(\u_cpu.rf_ram.memory[61][4] ),
    .A2(_03413_),
    .ZN(_03418_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08158_ (.A1(_03417_),
    .A2(_03407_),
    .B(_03418_),
    .ZN(_00347_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08159_ (.I(_03080_),
    .Z(_03419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08160_ (.A1(\u_cpu.rf_ram.memory[61][5] ),
    .A2(_03413_),
    .ZN(_03420_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08161_ (.A1(_03419_),
    .A2(_03408_),
    .B(_03420_),
    .ZN(_00348_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08162_ (.I(_03083_),
    .Z(_03421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08163_ (.A1(\u_cpu.rf_ram.memory[61][6] ),
    .A2(_03413_),
    .ZN(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08164_ (.A1(_03421_),
    .A2(_03408_),
    .B(_03422_),
    .ZN(_00349_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08165_ (.I(_03086_),
    .Z(_03423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08166_ (.A1(\u_cpu.rf_ram.memory[61][7] ),
    .A2(_03406_),
    .ZN(_03424_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08167_ (.A1(_03423_),
    .A2(_03408_),
    .B(_03424_),
    .ZN(_00350_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08168_ (.I(_03004_),
    .Z(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08169_ (.A1(_02981_),
    .A2(_03425_),
    .ZN(_03426_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08170_ (.I(_03426_),
    .Z(_03427_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08171_ (.I(_03426_),
    .Z(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08172_ (.A1(\u_cpu.rf_ram.memory[60][0] ),
    .A2(_03428_),
    .ZN(_03429_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08173_ (.A1(_03405_),
    .A2(_03427_),
    .B(_03429_),
    .ZN(_00351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08174_ (.A1(\u_cpu.rf_ram.memory[60][1] ),
    .A2(_03428_),
    .ZN(_03430_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08175_ (.A1(_03410_),
    .A2(_03427_),
    .B(_03430_),
    .ZN(_00352_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08176_ (.I(_03426_),
    .Z(_03431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08177_ (.A1(\u_cpu.rf_ram.memory[60][2] ),
    .A2(_03431_),
    .ZN(_03432_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08178_ (.A1(_03412_),
    .A2(_03427_),
    .B(_03432_),
    .ZN(_00353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08179_ (.A1(\u_cpu.rf_ram.memory[60][3] ),
    .A2(_03431_),
    .ZN(_03433_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08180_ (.A1(_03415_),
    .A2(_03427_),
    .B(_03433_),
    .ZN(_00354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08181_ (.A1(\u_cpu.rf_ram.memory[60][4] ),
    .A2(_03431_),
    .ZN(_03434_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08182_ (.A1(_03417_),
    .A2(_03427_),
    .B(_03434_),
    .ZN(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08183_ (.A1(\u_cpu.rf_ram.memory[60][5] ),
    .A2(_03431_),
    .ZN(_03435_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08184_ (.A1(_03419_),
    .A2(_03428_),
    .B(_03435_),
    .ZN(_00356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08185_ (.A1(\u_cpu.rf_ram.memory[60][6] ),
    .A2(_03431_),
    .ZN(_03436_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08186_ (.A1(_03421_),
    .A2(_03428_),
    .B(_03436_),
    .ZN(_00357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08187_ (.A1(\u_cpu.rf_ram.memory[60][7] ),
    .A2(_03426_),
    .ZN(_03437_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08188_ (.A1(_03423_),
    .A2(_03428_),
    .B(_03437_),
    .ZN(_00358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08189_ (.A1(_03367_),
    .A2(_03310_),
    .ZN(_03438_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08190_ (.I(_03438_),
    .Z(_03439_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08191_ (.I(_03438_),
    .Z(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08192_ (.A1(\u_cpu.rf_ram.memory[19][0] ),
    .A2(_03440_),
    .ZN(_03441_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08193_ (.A1(_03405_),
    .A2(_03439_),
    .B(_03441_),
    .ZN(_00359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08194_ (.A1(\u_cpu.rf_ram.memory[19][1] ),
    .A2(_03440_),
    .ZN(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08195_ (.A1(_03410_),
    .A2(_03439_),
    .B(_03442_),
    .ZN(_00360_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08196_ (.I(_03438_),
    .Z(_03443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08197_ (.A1(\u_cpu.rf_ram.memory[19][2] ),
    .A2(_03443_),
    .ZN(_03444_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08198_ (.A1(_03412_),
    .A2(_03439_),
    .B(_03444_),
    .ZN(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08199_ (.A1(\u_cpu.rf_ram.memory[19][3] ),
    .A2(_03443_),
    .ZN(_03445_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08200_ (.A1(_03415_),
    .A2(_03439_),
    .B(_03445_),
    .ZN(_00362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08201_ (.A1(\u_cpu.rf_ram.memory[19][4] ),
    .A2(_03443_),
    .ZN(_03446_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08202_ (.A1(_03417_),
    .A2(_03439_),
    .B(_03446_),
    .ZN(_00363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08203_ (.A1(\u_cpu.rf_ram.memory[19][5] ),
    .A2(_03443_),
    .ZN(_03447_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08204_ (.A1(_03419_),
    .A2(_03440_),
    .B(_03447_),
    .ZN(_00364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08205_ (.A1(\u_cpu.rf_ram.memory[19][6] ),
    .A2(_03443_),
    .ZN(_03448_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08206_ (.A1(_03421_),
    .A2(_03440_),
    .B(_03448_),
    .ZN(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08207_ (.A1(\u_cpu.rf_ram.memory[19][7] ),
    .A2(_03438_),
    .ZN(_03449_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08208_ (.A1(_03423_),
    .A2(_03440_),
    .B(_03449_),
    .ZN(_00366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08209_ (.A1(_02786_),
    .A2(_02850_),
    .ZN(_03450_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08210_ (.I(_03450_),
    .Z(_03451_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08211_ (.I0(_02846_),
    .I1(\u_cpu.rf_ram.memory[5][0] ),
    .S(_03451_),
    .Z(_03452_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08212_ (.I(_03452_),
    .Z(_00367_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08213_ (.I0(_02855_),
    .I1(\u_cpu.rf_ram.memory[5][1] ),
    .S(_03451_),
    .Z(_03453_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08214_ (.I(_03453_),
    .Z(_00368_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08215_ (.I0(_02858_),
    .I1(\u_cpu.rf_ram.memory[5][2] ),
    .S(_03451_),
    .Z(_03454_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08216_ (.I(_03454_),
    .Z(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08217_ (.I0(_02861_),
    .I1(\u_cpu.rf_ram.memory[5][3] ),
    .S(_03451_),
    .Z(_03455_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08218_ (.I(_03455_),
    .Z(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08219_ (.I0(_02864_),
    .I1(\u_cpu.rf_ram.memory[5][4] ),
    .S(_03451_),
    .Z(_03456_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08220_ (.I(_03456_),
    .Z(_00371_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08221_ (.I0(_02867_),
    .I1(\u_cpu.rf_ram.memory[5][5] ),
    .S(_03450_),
    .Z(_03457_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08222_ (.I(_03457_),
    .Z(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08223_ (.I0(_02870_),
    .I1(\u_cpu.rf_ram.memory[5][6] ),
    .S(_03450_),
    .Z(_03458_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08224_ (.I(_03458_),
    .Z(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08225_ (.I0(_02873_),
    .I1(\u_cpu.rf_ram.memory[5][7] ),
    .S(_03450_),
    .Z(_03459_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08226_ (.I(_03459_),
    .Z(_00374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08227_ (.A1(_02937_),
    .A2(_03425_),
    .ZN(_03460_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08228_ (.I(_03460_),
    .Z(_03461_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08229_ (.I(_03460_),
    .Z(_03462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08230_ (.A1(\u_cpu.rf_ram.memory[58][0] ),
    .A2(_03462_),
    .ZN(_03463_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08231_ (.A1(_03405_),
    .A2(_03461_),
    .B(_03463_),
    .ZN(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08232_ (.A1(\u_cpu.rf_ram.memory[58][1] ),
    .A2(_03462_),
    .ZN(_03464_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08233_ (.A1(_03410_),
    .A2(_03461_),
    .B(_03464_),
    .ZN(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08234_ (.I(_03460_),
    .Z(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08235_ (.A1(\u_cpu.rf_ram.memory[58][2] ),
    .A2(_03465_),
    .ZN(_03466_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08236_ (.A1(_03412_),
    .A2(_03461_),
    .B(_03466_),
    .ZN(_00377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08237_ (.A1(\u_cpu.rf_ram.memory[58][3] ),
    .A2(_03465_),
    .ZN(_03467_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08238_ (.A1(_03415_),
    .A2(_03461_),
    .B(_03467_),
    .ZN(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08239_ (.A1(\u_cpu.rf_ram.memory[58][4] ),
    .A2(_03465_),
    .ZN(_03468_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08240_ (.A1(_03417_),
    .A2(_03461_),
    .B(_03468_),
    .ZN(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08241_ (.A1(\u_cpu.rf_ram.memory[58][5] ),
    .A2(_03465_),
    .ZN(_03469_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08242_ (.A1(_03419_),
    .A2(_03462_),
    .B(_03469_),
    .ZN(_00380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08243_ (.A1(\u_cpu.rf_ram.memory[58][6] ),
    .A2(_03465_),
    .ZN(_03470_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08244_ (.A1(_03421_),
    .A2(_03462_),
    .B(_03470_),
    .ZN(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08245_ (.A1(\u_cpu.rf_ram.memory[58][7] ),
    .A2(_03460_),
    .ZN(_03471_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08246_ (.A1(_03423_),
    .A2(_03462_),
    .B(_03471_),
    .ZN(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08247_ (.A1(_03380_),
    .A2(_03020_),
    .ZN(_03472_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08248_ (.I(_03472_),
    .Z(_03473_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08249_ (.I(_03472_),
    .Z(_03474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08250_ (.A1(\u_cpu.rf_ram.memory[57][0] ),
    .A2(_03474_),
    .ZN(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08251_ (.A1(_03405_),
    .A2(_03473_),
    .B(_03475_),
    .ZN(_00383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08252_ (.A1(\u_cpu.rf_ram.memory[57][1] ),
    .A2(_03474_),
    .ZN(_03476_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08253_ (.A1(_03410_),
    .A2(_03473_),
    .B(_03476_),
    .ZN(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08254_ (.I(_03472_),
    .Z(_03477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08255_ (.A1(\u_cpu.rf_ram.memory[57][2] ),
    .A2(_03477_),
    .ZN(_03478_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08256_ (.A1(_03412_),
    .A2(_03473_),
    .B(_03478_),
    .ZN(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08257_ (.A1(\u_cpu.rf_ram.memory[57][3] ),
    .A2(_03477_),
    .ZN(_03479_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08258_ (.A1(_03415_),
    .A2(_03473_),
    .B(_03479_),
    .ZN(_00386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08259_ (.A1(\u_cpu.rf_ram.memory[57][4] ),
    .A2(_03477_),
    .ZN(_03480_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08260_ (.A1(_03417_),
    .A2(_03473_),
    .B(_03480_),
    .ZN(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08261_ (.A1(\u_cpu.rf_ram.memory[57][5] ),
    .A2(_03477_),
    .ZN(_03481_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08262_ (.A1(_03419_),
    .A2(_03474_),
    .B(_03481_),
    .ZN(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08263_ (.A1(\u_cpu.rf_ram.memory[57][6] ),
    .A2(_03477_),
    .ZN(_03482_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08264_ (.A1(_03421_),
    .A2(_03474_),
    .B(_03482_),
    .ZN(_00389_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08265_ (.A1(\u_cpu.rf_ram.memory[57][7] ),
    .A2(_03472_),
    .ZN(_03483_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08266_ (.A1(_03423_),
    .A2(_03474_),
    .B(_03483_),
    .ZN(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08267_ (.I(_02738_),
    .Z(_03484_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08268_ (.I(_03484_),
    .Z(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08269_ (.A1(_03380_),
    .A2(_03166_),
    .ZN(_03486_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08270_ (.I(_03486_),
    .Z(_03487_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08271_ (.I(_03486_),
    .Z(_03488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08272_ (.A1(\u_cpu.rf_ram.memory[56][0] ),
    .A2(_03488_),
    .ZN(_03489_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08273_ (.A1(_03485_),
    .A2(_03487_),
    .B(_03489_),
    .ZN(_00391_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08274_ (.I(_02744_),
    .Z(_03490_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08275_ (.I(_03490_),
    .Z(_03491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08276_ (.A1(\u_cpu.rf_ram.memory[56][1] ),
    .A2(_03488_),
    .ZN(_03492_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08277_ (.A1(_03491_),
    .A2(_03487_),
    .B(_03492_),
    .ZN(_00392_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08278_ (.I(_02750_),
    .Z(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08279_ (.I(_03493_),
    .Z(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08280_ (.I(_03486_),
    .Z(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08281_ (.A1(\u_cpu.rf_ram.memory[56][2] ),
    .A2(_03495_),
    .ZN(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08282_ (.A1(_03494_),
    .A2(_03487_),
    .B(_03496_),
    .ZN(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08283_ (.I(_02756_),
    .Z(_03497_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08284_ (.I(_03497_),
    .Z(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08285_ (.A1(\u_cpu.rf_ram.memory[56][3] ),
    .A2(_03495_),
    .ZN(_03499_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08286_ (.A1(_03498_),
    .A2(_03487_),
    .B(_03499_),
    .ZN(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08287_ (.I(_02761_),
    .Z(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08288_ (.I(_03500_),
    .Z(_03501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08289_ (.A1(\u_cpu.rf_ram.memory[56][4] ),
    .A2(_03495_),
    .ZN(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08290_ (.A1(_03501_),
    .A2(_03487_),
    .B(_03502_),
    .ZN(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08291_ (.I(_02766_),
    .Z(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08292_ (.I(_03503_),
    .Z(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08293_ (.A1(\u_cpu.rf_ram.memory[56][5] ),
    .A2(_03495_),
    .ZN(_03505_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08294_ (.A1(_03504_),
    .A2(_03488_),
    .B(_03505_),
    .ZN(_00396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08295_ (.I(_02771_),
    .Z(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08296_ (.I(_03506_),
    .Z(_03507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08297_ (.A1(\u_cpu.rf_ram.memory[56][6] ),
    .A2(_03495_),
    .ZN(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08298_ (.A1(_03507_),
    .A2(_03488_),
    .B(_03508_),
    .ZN(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08299_ (.I(_02776_),
    .Z(_03509_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08300_ (.I(_03509_),
    .Z(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08301_ (.A1(\u_cpu.rf_ram.memory[56][7] ),
    .A2(_03486_),
    .ZN(_03511_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08302_ (.A1(_03510_),
    .A2(_03488_),
    .B(_03511_),
    .ZN(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08303_ (.A1(_02877_),
    .A2(_03425_),
    .ZN(_03512_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08304_ (.I(_03512_),
    .Z(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08305_ (.I(_03512_),
    .Z(_03514_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08306_ (.A1(\u_cpu.rf_ram.memory[55][0] ),
    .A2(_03514_),
    .ZN(_03515_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08307_ (.A1(_03485_),
    .A2(_03513_),
    .B(_03515_),
    .ZN(_00399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08308_ (.A1(\u_cpu.rf_ram.memory[55][1] ),
    .A2(_03514_),
    .ZN(_03516_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08309_ (.A1(_03491_),
    .A2(_03513_),
    .B(_03516_),
    .ZN(_00400_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08310_ (.I(_03512_),
    .Z(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08311_ (.A1(\u_cpu.rf_ram.memory[55][2] ),
    .A2(_03517_),
    .ZN(_03518_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08312_ (.A1(_03494_),
    .A2(_03513_),
    .B(_03518_),
    .ZN(_00401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08313_ (.A1(\u_cpu.rf_ram.memory[55][3] ),
    .A2(_03517_),
    .ZN(_03519_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08314_ (.A1(_03498_),
    .A2(_03513_),
    .B(_03519_),
    .ZN(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08315_ (.A1(\u_cpu.rf_ram.memory[55][4] ),
    .A2(_03517_),
    .ZN(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08316_ (.A1(_03501_),
    .A2(_03513_),
    .B(_03520_),
    .ZN(_00403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08317_ (.A1(\u_cpu.rf_ram.memory[55][5] ),
    .A2(_03517_),
    .ZN(_03521_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08318_ (.A1(_03504_),
    .A2(_03514_),
    .B(_03521_),
    .ZN(_00404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08319_ (.A1(\u_cpu.rf_ram.memory[55][6] ),
    .A2(_03517_),
    .ZN(_03522_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08320_ (.A1(_03507_),
    .A2(_03514_),
    .B(_03522_),
    .ZN(_00405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08321_ (.A1(\u_cpu.rf_ram.memory[55][7] ),
    .A2(_03512_),
    .ZN(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08322_ (.A1(_03510_),
    .A2(_03514_),
    .B(_03523_),
    .ZN(_00406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08323_ (.A1(_03380_),
    .A2(_03287_),
    .ZN(_03524_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08324_ (.I(_03524_),
    .Z(_03525_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08325_ (.I(_03524_),
    .Z(_03526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08326_ (.A1(\u_cpu.rf_ram.memory[54][0] ),
    .A2(_03526_),
    .ZN(_03527_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08327_ (.A1(_03485_),
    .A2(_03525_),
    .B(_03527_),
    .ZN(_00407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08328_ (.A1(\u_cpu.rf_ram.memory[54][1] ),
    .A2(_03526_),
    .ZN(_03528_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08329_ (.A1(_03491_),
    .A2(_03525_),
    .B(_03528_),
    .ZN(_00408_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08330_ (.I(_03524_),
    .Z(_03529_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08331_ (.A1(\u_cpu.rf_ram.memory[54][2] ),
    .A2(_03529_),
    .ZN(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08332_ (.A1(_03494_),
    .A2(_03525_),
    .B(_03530_),
    .ZN(_00409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08333_ (.A1(\u_cpu.rf_ram.memory[54][3] ),
    .A2(_03529_),
    .ZN(_03531_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08334_ (.A1(_03498_),
    .A2(_03525_),
    .B(_03531_),
    .ZN(_00410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08335_ (.A1(\u_cpu.rf_ram.memory[54][4] ),
    .A2(_03529_),
    .ZN(_03532_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08336_ (.A1(_03501_),
    .A2(_03525_),
    .B(_03532_),
    .ZN(_00411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08337_ (.A1(\u_cpu.rf_ram.memory[54][5] ),
    .A2(_03529_),
    .ZN(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08338_ (.A1(_03504_),
    .A2(_03526_),
    .B(_03533_),
    .ZN(_00412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08339_ (.A1(\u_cpu.rf_ram.memory[54][6] ),
    .A2(_03529_),
    .ZN(_03534_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08340_ (.A1(_03507_),
    .A2(_03526_),
    .B(_03534_),
    .ZN(_00413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08341_ (.A1(\u_cpu.rf_ram.memory[54][7] ),
    .A2(_03524_),
    .ZN(_03535_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08342_ (.A1(_03510_),
    .A2(_03526_),
    .B(_03535_),
    .ZN(_00414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08343_ (.A1(_02786_),
    .A2(_03425_),
    .ZN(_03536_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08344_ (.I(_03536_),
    .Z(_03537_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08345_ (.I(_03536_),
    .Z(_03538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08346_ (.A1(\u_cpu.rf_ram.memory[53][0] ),
    .A2(_03538_),
    .ZN(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08347_ (.A1(_03485_),
    .A2(_03537_),
    .B(_03539_),
    .ZN(_00415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08348_ (.A1(\u_cpu.rf_ram.memory[53][1] ),
    .A2(_03538_),
    .ZN(_03540_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08349_ (.A1(_03491_),
    .A2(_03537_),
    .B(_03540_),
    .ZN(_00416_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08350_ (.I(_03536_),
    .Z(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08351_ (.A1(\u_cpu.rf_ram.memory[53][2] ),
    .A2(_03541_),
    .ZN(_03542_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08352_ (.A1(_03494_),
    .A2(_03537_),
    .B(_03542_),
    .ZN(_00417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08353_ (.A1(\u_cpu.rf_ram.memory[53][3] ),
    .A2(_03541_),
    .ZN(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08354_ (.A1(_03498_),
    .A2(_03537_),
    .B(_03543_),
    .ZN(_00418_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08355_ (.A1(\u_cpu.rf_ram.memory[53][4] ),
    .A2(_03541_),
    .ZN(_03544_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08356_ (.A1(_03501_),
    .A2(_03537_),
    .B(_03544_),
    .ZN(_00419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08357_ (.A1(\u_cpu.rf_ram.memory[53][5] ),
    .A2(_03541_),
    .ZN(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08358_ (.A1(_03504_),
    .A2(_03538_),
    .B(_03545_),
    .ZN(_00420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08359_ (.A1(\u_cpu.rf_ram.memory[53][6] ),
    .A2(_03541_),
    .ZN(_03546_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08360_ (.A1(_03507_),
    .A2(_03538_),
    .B(_03546_),
    .ZN(_00421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08361_ (.A1(\u_cpu.rf_ram.memory[53][7] ),
    .A2(_03536_),
    .ZN(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08362_ (.A1(_03510_),
    .A2(_03538_),
    .B(_03547_),
    .ZN(_00422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08363_ (.A1(_02831_),
    .A2(_03425_),
    .ZN(_03548_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08364_ (.I(_03548_),
    .Z(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08365_ (.I(_03548_),
    .Z(_03550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08366_ (.A1(\u_cpu.rf_ram.memory[52][0] ),
    .A2(_03550_),
    .ZN(_03551_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08367_ (.A1(_03485_),
    .A2(_03549_),
    .B(_03551_),
    .ZN(_00423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08368_ (.A1(\u_cpu.rf_ram.memory[52][1] ),
    .A2(_03550_),
    .ZN(_03552_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08369_ (.A1(_03491_),
    .A2(_03549_),
    .B(_03552_),
    .ZN(_00424_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08370_ (.I(_03548_),
    .Z(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08371_ (.A1(\u_cpu.rf_ram.memory[52][2] ),
    .A2(_03553_),
    .ZN(_03554_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08372_ (.A1(_03494_),
    .A2(_03549_),
    .B(_03554_),
    .ZN(_00425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08373_ (.A1(\u_cpu.rf_ram.memory[52][3] ),
    .A2(_03553_),
    .ZN(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08374_ (.A1(_03498_),
    .A2(_03549_),
    .B(_03555_),
    .ZN(_00426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08375_ (.A1(\u_cpu.rf_ram.memory[52][4] ),
    .A2(_03553_),
    .ZN(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08376_ (.A1(_03501_),
    .A2(_03549_),
    .B(_03556_),
    .ZN(_00427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08377_ (.A1(\u_cpu.rf_ram.memory[52][5] ),
    .A2(_03553_),
    .ZN(_03557_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08378_ (.A1(_03504_),
    .A2(_03550_),
    .B(_03557_),
    .ZN(_00428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08379_ (.A1(\u_cpu.rf_ram.memory[52][6] ),
    .A2(_03553_),
    .ZN(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08380_ (.A1(_03507_),
    .A2(_03550_),
    .B(_03558_),
    .ZN(_00429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08381_ (.A1(\u_cpu.rf_ram.memory[52][7] ),
    .A2(_03548_),
    .ZN(_03559_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08382_ (.A1(_03510_),
    .A2(_03550_),
    .B(_03559_),
    .ZN(_00430_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08383_ (.I(_02845_),
    .Z(_03560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08384_ (.A1(_03285_),
    .A2(_03020_),
    .ZN(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08385_ (.I(_03561_),
    .Z(_03562_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08386_ (.I0(_03560_),
    .I1(\u_cpu.rf_ram.memory[9][0] ),
    .S(_03562_),
    .Z(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08387_ (.I(_03563_),
    .Z(_00431_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08388_ (.I(_02854_),
    .Z(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08389_ (.I0(_03564_),
    .I1(\u_cpu.rf_ram.memory[9][1] ),
    .S(_03562_),
    .Z(_03565_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08390_ (.I(_03565_),
    .Z(_00432_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08391_ (.I(_02857_),
    .Z(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08392_ (.I0(_03566_),
    .I1(\u_cpu.rf_ram.memory[9][2] ),
    .S(_03562_),
    .Z(_03567_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08393_ (.I(_03567_),
    .Z(_00433_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08394_ (.I(_02860_),
    .Z(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08395_ (.I0(_03568_),
    .I1(\u_cpu.rf_ram.memory[9][3] ),
    .S(_03562_),
    .Z(_03569_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08396_ (.I(_03569_),
    .Z(_00434_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08397_ (.I(_02863_),
    .Z(_03570_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08398_ (.I0(_03570_),
    .I1(\u_cpu.rf_ram.memory[9][4] ),
    .S(_03562_),
    .Z(_03571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08399_ (.I(_03571_),
    .Z(_00435_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08400_ (.I(_02866_),
    .Z(_03572_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08401_ (.I0(_03572_),
    .I1(\u_cpu.rf_ram.memory[9][5] ),
    .S(_03561_),
    .Z(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08402_ (.I(_03573_),
    .Z(_00436_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08403_ (.I(_02869_),
    .Z(_03574_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08404_ (.I0(_03574_),
    .I1(\u_cpu.rf_ram.memory[9][6] ),
    .S(_03561_),
    .Z(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08405_ (.I(_03575_),
    .Z(_00437_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08406_ (.I(_02872_),
    .Z(_03576_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08407_ (.I0(_03576_),
    .I1(\u_cpu.rf_ram.memory[9][7] ),
    .S(_03561_),
    .Z(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08408_ (.I(_03577_),
    .Z(_00438_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08409_ (.A1(_03285_),
    .A2(_03062_),
    .ZN(_03578_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08410_ (.I(_03578_),
    .Z(_03579_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08411_ (.I0(_03560_),
    .I1(\u_cpu.rf_ram.memory[15][0] ),
    .S(_03579_),
    .Z(_03580_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08412_ (.I(_03580_),
    .Z(_00439_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08413_ (.I0(_03564_),
    .I1(\u_cpu.rf_ram.memory[15][1] ),
    .S(_03579_),
    .Z(_03581_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08414_ (.I(_03581_),
    .Z(_00440_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08415_ (.I0(_03566_),
    .I1(\u_cpu.rf_ram.memory[15][2] ),
    .S(_03579_),
    .Z(_03582_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08416_ (.I(_03582_),
    .Z(_00441_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08417_ (.I0(_03568_),
    .I1(\u_cpu.rf_ram.memory[15][3] ),
    .S(_03579_),
    .Z(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08418_ (.I(_03583_),
    .Z(_00442_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08419_ (.I0(_03570_),
    .I1(\u_cpu.rf_ram.memory[15][4] ),
    .S(_03579_),
    .Z(_03584_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08420_ (.I(_03584_),
    .Z(_00443_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08421_ (.I0(_03572_),
    .I1(\u_cpu.rf_ram.memory[15][5] ),
    .S(_03578_),
    .Z(_03585_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08422_ (.I(_03585_),
    .Z(_00444_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08423_ (.I0(_03574_),
    .I1(\u_cpu.rf_ram.memory[15][6] ),
    .S(_03578_),
    .Z(_03586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08424_ (.I(_03586_),
    .Z(_00445_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08425_ (.I0(_03576_),
    .I1(\u_cpu.rf_ram.memory[15][7] ),
    .S(_03578_),
    .Z(_03587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08426_ (.I(_03587_),
    .Z(_00446_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08427_ (.I(_03484_),
    .Z(_03588_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08428_ (.A1(_02920_),
    .A2(_03202_),
    .ZN(_03589_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08429_ (.I(_03589_),
    .Z(_03590_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08430_ (.I(_03589_),
    .Z(_03591_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08431_ (.A1(\u_cpu.rf_ram.memory[142][0] ),
    .A2(_03591_),
    .ZN(_03592_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08432_ (.A1(_03588_),
    .A2(_03590_),
    .B(_03592_),
    .ZN(_00447_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08433_ (.I(_03490_),
    .Z(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08434_ (.A1(\u_cpu.rf_ram.memory[142][1] ),
    .A2(_03591_),
    .ZN(_03594_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08435_ (.A1(_03593_),
    .A2(_03590_),
    .B(_03594_),
    .ZN(_00448_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08436_ (.I(_03493_),
    .Z(_03595_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08437_ (.I(_03589_),
    .Z(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08438_ (.A1(\u_cpu.rf_ram.memory[142][2] ),
    .A2(_03596_),
    .ZN(_03597_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08439_ (.A1(_03595_),
    .A2(_03590_),
    .B(_03597_),
    .ZN(_00449_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08440_ (.I(_03497_),
    .Z(_03598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08441_ (.A1(\u_cpu.rf_ram.memory[142][3] ),
    .A2(_03596_),
    .ZN(_03599_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08442_ (.A1(_03598_),
    .A2(_03590_),
    .B(_03599_),
    .ZN(_00450_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08443_ (.I(_03500_),
    .Z(_03600_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08444_ (.A1(\u_cpu.rf_ram.memory[142][4] ),
    .A2(_03596_),
    .ZN(_03601_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08445_ (.A1(_03600_),
    .A2(_03590_),
    .B(_03601_),
    .ZN(_00451_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08446_ (.I(_03503_),
    .Z(_03602_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08447_ (.A1(\u_cpu.rf_ram.memory[142][5] ),
    .A2(_03596_),
    .ZN(_03603_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08448_ (.A1(_03602_),
    .A2(_03591_),
    .B(_03603_),
    .ZN(_00452_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08449_ (.I(_03506_),
    .Z(_03604_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08450_ (.A1(\u_cpu.rf_ram.memory[142][6] ),
    .A2(_03596_),
    .ZN(_03605_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08451_ (.A1(_03604_),
    .A2(_03591_),
    .B(_03605_),
    .ZN(_00453_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08452_ (.I(_03509_),
    .Z(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08453_ (.A1(\u_cpu.rf_ram.memory[142][7] ),
    .A2(_03589_),
    .ZN(_03607_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08454_ (.A1(_03606_),
    .A2(_03591_),
    .B(_03607_),
    .ZN(_00454_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08455_ (.A1(_02966_),
    .A2(_03202_),
    .ZN(_03608_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08456_ (.I(_03608_),
    .Z(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08457_ (.I(_03608_),
    .Z(_03610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08458_ (.A1(\u_cpu.rf_ram.memory[141][0] ),
    .A2(_03610_),
    .ZN(_03611_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08459_ (.A1(_03588_),
    .A2(_03609_),
    .B(_03611_),
    .ZN(_00455_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08460_ (.A1(\u_cpu.rf_ram.memory[141][1] ),
    .A2(_03610_),
    .ZN(_03612_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08461_ (.A1(_03593_),
    .A2(_03609_),
    .B(_03612_),
    .ZN(_00456_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08462_ (.I(_03608_),
    .Z(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08463_ (.A1(\u_cpu.rf_ram.memory[141][2] ),
    .A2(_03613_),
    .ZN(_03614_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08464_ (.A1(_03595_),
    .A2(_03609_),
    .B(_03614_),
    .ZN(_00457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08465_ (.A1(\u_cpu.rf_ram.memory[141][3] ),
    .A2(_03613_),
    .ZN(_03615_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08466_ (.A1(_03598_),
    .A2(_03609_),
    .B(_03615_),
    .ZN(_00458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08467_ (.A1(\u_cpu.rf_ram.memory[141][4] ),
    .A2(_03613_),
    .ZN(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08468_ (.A1(_03600_),
    .A2(_03609_),
    .B(_03616_),
    .ZN(_00459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08469_ (.A1(\u_cpu.rf_ram.memory[141][5] ),
    .A2(_03613_),
    .ZN(_03617_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08470_ (.A1(_03602_),
    .A2(_03610_),
    .B(_03617_),
    .ZN(_00460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08471_ (.A1(\u_cpu.rf_ram.memory[141][6] ),
    .A2(_03613_),
    .ZN(_03618_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08472_ (.A1(_03604_),
    .A2(_03610_),
    .B(_03618_),
    .ZN(_00461_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08473_ (.A1(\u_cpu.rf_ram.memory[141][7] ),
    .A2(_03608_),
    .ZN(_03619_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08474_ (.A1(_03606_),
    .A2(_03610_),
    .B(_03619_),
    .ZN(_00462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08475_ (.A1(_02981_),
    .A2(_03202_),
    .ZN(_03620_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08476_ (.I(_03620_),
    .Z(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08477_ (.I(_03620_),
    .Z(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08478_ (.A1(\u_cpu.rf_ram.memory[140][0] ),
    .A2(_03622_),
    .ZN(_03623_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08479_ (.A1(_03588_),
    .A2(_03621_),
    .B(_03623_),
    .ZN(_00463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08480_ (.A1(\u_cpu.rf_ram.memory[140][1] ),
    .A2(_03622_),
    .ZN(_03624_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08481_ (.A1(_03593_),
    .A2(_03621_),
    .B(_03624_),
    .ZN(_00464_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08482_ (.I(_03620_),
    .Z(_03625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08483_ (.A1(\u_cpu.rf_ram.memory[140][2] ),
    .A2(_03625_),
    .ZN(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08484_ (.A1(_03595_),
    .A2(_03621_),
    .B(_03626_),
    .ZN(_00465_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08485_ (.A1(\u_cpu.rf_ram.memory[140][3] ),
    .A2(_03625_),
    .ZN(_03627_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08486_ (.A1(_03598_),
    .A2(_03621_),
    .B(_03627_),
    .ZN(_00466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08487_ (.A1(\u_cpu.rf_ram.memory[140][4] ),
    .A2(_03625_),
    .ZN(_03628_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08488_ (.A1(_03600_),
    .A2(_03621_),
    .B(_03628_),
    .ZN(_00467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08489_ (.A1(\u_cpu.rf_ram.memory[140][5] ),
    .A2(_03625_),
    .ZN(_03629_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08490_ (.A1(_03602_),
    .A2(_03622_),
    .B(_03629_),
    .ZN(_00468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08491_ (.A1(\u_cpu.rf_ram.memory[140][6] ),
    .A2(_03625_),
    .ZN(_03630_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08492_ (.A1(_03604_),
    .A2(_03622_),
    .B(_03630_),
    .ZN(_00469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08493_ (.A1(\u_cpu.rf_ram.memory[140][7] ),
    .A2(_03620_),
    .ZN(_03631_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08494_ (.A1(_03606_),
    .A2(_03622_),
    .B(_03631_),
    .ZN(_00470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08495_ (.A1(_03285_),
    .A2(_02967_),
    .ZN(_03632_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08496_ (.I(_03632_),
    .Z(_03633_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08497_ (.I0(_03560_),
    .I1(\u_cpu.rf_ram.memory[13][0] ),
    .S(_03633_),
    .Z(_03634_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08498_ (.I(_03634_),
    .Z(_00471_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08499_ (.I0(_03564_),
    .I1(\u_cpu.rf_ram.memory[13][1] ),
    .S(_03633_),
    .Z(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08500_ (.I(_03635_),
    .Z(_00472_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08501_ (.I0(_03566_),
    .I1(\u_cpu.rf_ram.memory[13][2] ),
    .S(_03633_),
    .Z(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08502_ (.I(_03636_),
    .Z(_00473_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08503_ (.I0(_03568_),
    .I1(\u_cpu.rf_ram.memory[13][3] ),
    .S(_03633_),
    .Z(_03637_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08504_ (.I(_03637_),
    .Z(_00474_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08505_ (.I0(_03570_),
    .I1(\u_cpu.rf_ram.memory[13][4] ),
    .S(_03633_),
    .Z(_03638_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08506_ (.I(_03638_),
    .Z(_00475_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08507_ (.I0(_03572_),
    .I1(\u_cpu.rf_ram.memory[13][5] ),
    .S(_03632_),
    .Z(_03639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08508_ (.I(_03639_),
    .Z(_00476_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08509_ (.I0(_03574_),
    .I1(\u_cpu.rf_ram.memory[13][6] ),
    .S(_03632_),
    .Z(_03640_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08510_ (.I(_03640_),
    .Z(_00477_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08511_ (.I0(_03576_),
    .I1(\u_cpu.rf_ram.memory[13][7] ),
    .S(_03632_),
    .Z(_03641_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08512_ (.I(_03641_),
    .Z(_00478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08513_ (.A1(_03272_),
    .A2(_03166_),
    .ZN(_03642_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08514_ (.I(_03642_),
    .Z(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08515_ (.I(_03642_),
    .Z(_03644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08516_ (.A1(\u_cpu.rf_ram.memory[72][0] ),
    .A2(_03644_),
    .ZN(_03645_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08517_ (.A1(_03588_),
    .A2(_03643_),
    .B(_03645_),
    .ZN(_00479_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08518_ (.A1(\u_cpu.rf_ram.memory[72][1] ),
    .A2(_03644_),
    .ZN(_03646_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08519_ (.A1(_03593_),
    .A2(_03643_),
    .B(_03646_),
    .ZN(_00480_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08520_ (.I(_03642_),
    .Z(_03647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08521_ (.A1(\u_cpu.rf_ram.memory[72][2] ),
    .A2(_03647_),
    .ZN(_03648_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08522_ (.A1(_03595_),
    .A2(_03643_),
    .B(_03648_),
    .ZN(_00481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08523_ (.A1(\u_cpu.rf_ram.memory[72][3] ),
    .A2(_03647_),
    .ZN(_03649_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08524_ (.A1(_03598_),
    .A2(_03643_),
    .B(_03649_),
    .ZN(_00482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08525_ (.A1(\u_cpu.rf_ram.memory[72][4] ),
    .A2(_03647_),
    .ZN(_03650_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08526_ (.A1(_03600_),
    .A2(_03643_),
    .B(_03650_),
    .ZN(_00483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08527_ (.A1(\u_cpu.rf_ram.memory[72][5] ),
    .A2(_03647_),
    .ZN(_03651_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08528_ (.A1(_03602_),
    .A2(_03644_),
    .B(_03651_),
    .ZN(_00484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08529_ (.A1(\u_cpu.rf_ram.memory[72][6] ),
    .A2(_03647_),
    .ZN(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08530_ (.A1(_03604_),
    .A2(_03644_),
    .B(_03652_),
    .ZN(_00485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08531_ (.A1(\u_cpu.rf_ram.memory[72][7] ),
    .A2(_03642_),
    .ZN(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08532_ (.A1(_03606_),
    .A2(_03644_),
    .B(_03653_),
    .ZN(_00486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08533_ (.A1(_03272_),
    .A2(_03020_),
    .ZN(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08534_ (.I(_03654_),
    .Z(_03655_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08535_ (.I(_03654_),
    .Z(_03656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08536_ (.A1(\u_cpu.rf_ram.memory[73][0] ),
    .A2(_03656_),
    .ZN(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08537_ (.A1(_03588_),
    .A2(_03655_),
    .B(_03657_),
    .ZN(_00487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08538_ (.A1(\u_cpu.rf_ram.memory[73][1] ),
    .A2(_03656_),
    .ZN(_03658_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08539_ (.A1(_03593_),
    .A2(_03655_),
    .B(_03658_),
    .ZN(_00488_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08540_ (.I(_03654_),
    .Z(_03659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08541_ (.A1(\u_cpu.rf_ram.memory[73][2] ),
    .A2(_03659_),
    .ZN(_03660_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08542_ (.A1(_03595_),
    .A2(_03655_),
    .B(_03660_),
    .ZN(_00489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08543_ (.A1(\u_cpu.rf_ram.memory[73][3] ),
    .A2(_03659_),
    .ZN(_03661_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08544_ (.A1(_03598_),
    .A2(_03655_),
    .B(_03661_),
    .ZN(_00490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08545_ (.A1(\u_cpu.rf_ram.memory[73][4] ),
    .A2(_03659_),
    .ZN(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08546_ (.A1(_03600_),
    .A2(_03655_),
    .B(_03662_),
    .ZN(_00491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08547_ (.A1(\u_cpu.rf_ram.memory[73][5] ),
    .A2(_03659_),
    .ZN(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08548_ (.A1(_03602_),
    .A2(_03656_),
    .B(_03663_),
    .ZN(_00492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08549_ (.A1(\u_cpu.rf_ram.memory[73][6] ),
    .A2(_03659_),
    .ZN(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08550_ (.A1(_03604_),
    .A2(_03656_),
    .B(_03664_),
    .ZN(_00493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08551_ (.A1(\u_cpu.rf_ram.memory[73][7] ),
    .A2(_03654_),
    .ZN(_03665_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08552_ (.A1(_03606_),
    .A2(_03656_),
    .B(_03665_),
    .ZN(_00494_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08553_ (.I(_03484_),
    .Z(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08554_ (.A1(_02876_),
    .A2(_03227_),
    .ZN(_03667_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08555_ (.I(_03667_),
    .Z(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08556_ (.I(_03667_),
    .Z(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08557_ (.A1(\u_cpu.rf_ram.memory[71][0] ),
    .A2(_03669_),
    .ZN(_03670_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08558_ (.A1(_03666_),
    .A2(_03668_),
    .B(_03670_),
    .ZN(_00495_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08559_ (.I(_03490_),
    .Z(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08560_ (.A1(\u_cpu.rf_ram.memory[71][1] ),
    .A2(_03669_),
    .ZN(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08561_ (.A1(_03671_),
    .A2(_03668_),
    .B(_03672_),
    .ZN(_00496_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08562_ (.I(_03493_),
    .Z(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08563_ (.I(_03667_),
    .Z(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08564_ (.A1(\u_cpu.rf_ram.memory[71][2] ),
    .A2(_03674_),
    .ZN(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08565_ (.A1(_03673_),
    .A2(_03668_),
    .B(_03675_),
    .ZN(_00497_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08566_ (.I(_03497_),
    .Z(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08567_ (.A1(\u_cpu.rf_ram.memory[71][3] ),
    .A2(_03674_),
    .ZN(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08568_ (.A1(_03676_),
    .A2(_03668_),
    .B(_03677_),
    .ZN(_00498_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08569_ (.I(_03500_),
    .Z(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08570_ (.A1(\u_cpu.rf_ram.memory[71][4] ),
    .A2(_03674_),
    .ZN(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08571_ (.A1(_03678_),
    .A2(_03668_),
    .B(_03679_),
    .ZN(_00499_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08572_ (.I(_03503_),
    .Z(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08573_ (.A1(\u_cpu.rf_ram.memory[71][5] ),
    .A2(_03674_),
    .ZN(_03681_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08574_ (.A1(_03680_),
    .A2(_03669_),
    .B(_03681_),
    .ZN(_00500_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08575_ (.I(_03506_),
    .Z(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08576_ (.A1(\u_cpu.rf_ram.memory[71][6] ),
    .A2(_03674_),
    .ZN(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08577_ (.A1(_03682_),
    .A2(_03669_),
    .B(_03683_),
    .ZN(_00501_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08578_ (.I(_03509_),
    .Z(_03684_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08579_ (.A1(\u_cpu.rf_ram.memory[71][7] ),
    .A2(_03667_),
    .ZN(_03685_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08580_ (.A1(_03684_),
    .A2(_03669_),
    .B(_03685_),
    .ZN(_00502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08581_ (.A1(_03272_),
    .A2(_03287_),
    .ZN(_03686_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08582_ (.I(_03686_),
    .Z(_03687_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08583_ (.I(_03686_),
    .Z(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08584_ (.A1(\u_cpu.rf_ram.memory[70][0] ),
    .A2(_03688_),
    .ZN(_03689_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08585_ (.A1(_03666_),
    .A2(_03687_),
    .B(_03689_),
    .ZN(_00503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08586_ (.A1(\u_cpu.rf_ram.memory[70][1] ),
    .A2(_03688_),
    .ZN(_03690_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08587_ (.A1(_03671_),
    .A2(_03687_),
    .B(_03690_),
    .ZN(_00504_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08588_ (.I(_03686_),
    .Z(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08589_ (.A1(\u_cpu.rf_ram.memory[70][2] ),
    .A2(_03691_),
    .ZN(_03692_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08590_ (.A1(_03673_),
    .A2(_03687_),
    .B(_03692_),
    .ZN(_00505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08591_ (.A1(\u_cpu.rf_ram.memory[70][3] ),
    .A2(_03691_),
    .ZN(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08592_ (.A1(_03676_),
    .A2(_03687_),
    .B(_03693_),
    .ZN(_00506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08593_ (.A1(\u_cpu.rf_ram.memory[70][4] ),
    .A2(_03691_),
    .ZN(_03694_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08594_ (.A1(_03678_),
    .A2(_03687_),
    .B(_03694_),
    .ZN(_00507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08595_ (.A1(\u_cpu.rf_ram.memory[70][5] ),
    .A2(_03691_),
    .ZN(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08596_ (.A1(_03680_),
    .A2(_03688_),
    .B(_03695_),
    .ZN(_00508_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08597_ (.A1(\u_cpu.rf_ram.memory[70][6] ),
    .A2(_03691_),
    .ZN(_03696_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08598_ (.A1(_03682_),
    .A2(_03688_),
    .B(_03696_),
    .ZN(_00509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08599_ (.A1(\u_cpu.rf_ram.memory[70][7] ),
    .A2(_03686_),
    .ZN(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08600_ (.A1(_03684_),
    .A2(_03688_),
    .B(_03697_),
    .ZN(_00510_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08601_ (.I(_03201_),
    .Z(_03698_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08602_ (.A1(_03061_),
    .A2(_03698_),
    .ZN(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08603_ (.I(_03699_),
    .Z(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08604_ (.I(_03699_),
    .Z(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08605_ (.A1(\u_cpu.rf_ram.memory[143][0] ),
    .A2(_03701_),
    .ZN(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08606_ (.A1(_03666_),
    .A2(_03700_),
    .B(_03702_),
    .ZN(_00511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08607_ (.A1(\u_cpu.rf_ram.memory[143][1] ),
    .A2(_03701_),
    .ZN(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08608_ (.A1(_03671_),
    .A2(_03700_),
    .B(_03703_),
    .ZN(_00512_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08609_ (.I(_03699_),
    .Z(_03704_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08610_ (.A1(\u_cpu.rf_ram.memory[143][2] ),
    .A2(_03704_),
    .ZN(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08611_ (.A1(_03673_),
    .A2(_03700_),
    .B(_03705_),
    .ZN(_00513_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08612_ (.A1(\u_cpu.rf_ram.memory[143][3] ),
    .A2(_03704_),
    .ZN(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08613_ (.A1(_03676_),
    .A2(_03700_),
    .B(_03706_),
    .ZN(_00514_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08614_ (.A1(\u_cpu.rf_ram.memory[143][4] ),
    .A2(_03704_),
    .ZN(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08615_ (.A1(_03678_),
    .A2(_03700_),
    .B(_03707_),
    .ZN(_00515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08616_ (.A1(\u_cpu.rf_ram.memory[143][5] ),
    .A2(_03704_),
    .ZN(_03708_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08617_ (.A1(_03680_),
    .A2(_03701_),
    .B(_03708_),
    .ZN(_00516_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08618_ (.A1(\u_cpu.rf_ram.memory[143][6] ),
    .A2(_03704_),
    .ZN(_03709_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08619_ (.A1(_03682_),
    .A2(_03701_),
    .B(_03709_),
    .ZN(_00517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08620_ (.A1(\u_cpu.rf_ram.memory[143][7] ),
    .A2(_03699_),
    .ZN(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08621_ (.A1(_03684_),
    .A2(_03701_),
    .B(_03710_),
    .ZN(_00518_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08622_ (.A1(_03285_),
    .A2(_02921_),
    .ZN(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08623_ (.I(_03711_),
    .Z(_03712_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08624_ (.I0(_03560_),
    .I1(\u_cpu.rf_ram.memory[14][0] ),
    .S(_03712_),
    .Z(_03713_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08625_ (.I(_03713_),
    .Z(_00519_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08626_ (.I0(_03564_),
    .I1(\u_cpu.rf_ram.memory[14][1] ),
    .S(_03712_),
    .Z(_03714_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08627_ (.I(_03714_),
    .Z(_00520_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08628_ (.I0(_03566_),
    .I1(\u_cpu.rf_ram.memory[14][2] ),
    .S(_03712_),
    .Z(_03715_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08629_ (.I(_03715_),
    .Z(_00521_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08630_ (.I0(_03568_),
    .I1(\u_cpu.rf_ram.memory[14][3] ),
    .S(_03712_),
    .Z(_03716_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08631_ (.I(_03716_),
    .Z(_00522_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08632_ (.I0(_03570_),
    .I1(\u_cpu.rf_ram.memory[14][4] ),
    .S(_03712_),
    .Z(_03717_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08633_ (.I(_03717_),
    .Z(_00523_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08634_ (.I0(_03572_),
    .I1(\u_cpu.rf_ram.memory[14][5] ),
    .S(_03711_),
    .Z(_03718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08635_ (.I(_03718_),
    .Z(_00524_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08636_ (.I0(_03574_),
    .I1(\u_cpu.rf_ram.memory[14][6] ),
    .S(_03711_),
    .Z(_03719_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08637_ (.I(_03719_),
    .Z(_00525_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08638_ (.I0(_03576_),
    .I1(\u_cpu.rf_ram.memory[14][7] ),
    .S(_03711_),
    .Z(_03720_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08639_ (.I(_03720_),
    .Z(_00526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08640_ (.A1(_02937_),
    .A2(_03698_),
    .ZN(_03721_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08641_ (.I(_03721_),
    .Z(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08642_ (.I(_03721_),
    .Z(_03723_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08643_ (.A1(\u_cpu.rf_ram.memory[138][0] ),
    .A2(_03723_),
    .ZN(_03724_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08644_ (.A1(_03666_),
    .A2(_03722_),
    .B(_03724_),
    .ZN(_00527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08645_ (.A1(\u_cpu.rf_ram.memory[138][1] ),
    .A2(_03723_),
    .ZN(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08646_ (.A1(_03671_),
    .A2(_03722_),
    .B(_03725_),
    .ZN(_00528_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08647_ (.I(_03721_),
    .Z(_03726_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08648_ (.A1(\u_cpu.rf_ram.memory[138][2] ),
    .A2(_03726_),
    .ZN(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08649_ (.A1(_03673_),
    .A2(_03722_),
    .B(_03727_),
    .ZN(_00529_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08650_ (.A1(\u_cpu.rf_ram.memory[138][3] ),
    .A2(_03726_),
    .ZN(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08651_ (.A1(_03676_),
    .A2(_03722_),
    .B(_03728_),
    .ZN(_00530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08652_ (.A1(\u_cpu.rf_ram.memory[138][4] ),
    .A2(_03726_),
    .ZN(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08653_ (.A1(_03678_),
    .A2(_03722_),
    .B(_03729_),
    .ZN(_00531_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08654_ (.A1(\u_cpu.rf_ram.memory[138][5] ),
    .A2(_03726_),
    .ZN(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08655_ (.A1(_03680_),
    .A2(_03723_),
    .B(_03730_),
    .ZN(_00532_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08656_ (.A1(\u_cpu.rf_ram.memory[138][6] ),
    .A2(_03726_),
    .ZN(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08657_ (.A1(_03682_),
    .A2(_03723_),
    .B(_03731_),
    .ZN(_00533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08658_ (.A1(\u_cpu.rf_ram.memory[138][7] ),
    .A2(_03721_),
    .ZN(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08659_ (.A1(_03684_),
    .A2(_03723_),
    .B(_03732_),
    .ZN(_00534_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08660_ (.A1(_02876_),
    .A2(_02940_),
    .ZN(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08661_ (.I(_03733_),
    .Z(_03734_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08662_ (.I(_03733_),
    .Z(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08663_ (.A1(\u_cpu.rf_ram.memory[39][0] ),
    .A2(_03735_),
    .ZN(_03736_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08664_ (.A1(_03666_),
    .A2(_03734_),
    .B(_03736_),
    .ZN(_00535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08665_ (.A1(\u_cpu.rf_ram.memory[39][1] ),
    .A2(_03735_),
    .ZN(_03737_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08666_ (.A1(_03671_),
    .A2(_03734_),
    .B(_03737_),
    .ZN(_00536_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08667_ (.I(_03733_),
    .Z(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08668_ (.A1(\u_cpu.rf_ram.memory[39][2] ),
    .A2(_03738_),
    .ZN(_03739_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08669_ (.A1(_03673_),
    .A2(_03734_),
    .B(_03739_),
    .ZN(_00537_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08670_ (.A1(\u_cpu.rf_ram.memory[39][3] ),
    .A2(_03738_),
    .ZN(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08671_ (.A1(_03676_),
    .A2(_03734_),
    .B(_03740_),
    .ZN(_00538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08672_ (.A1(\u_cpu.rf_ram.memory[39][4] ),
    .A2(_03738_),
    .ZN(_03741_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08673_ (.A1(_03678_),
    .A2(_03734_),
    .B(_03741_),
    .ZN(_00539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08674_ (.A1(\u_cpu.rf_ram.memory[39][5] ),
    .A2(_03738_),
    .ZN(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08675_ (.A1(_03680_),
    .A2(_03735_),
    .B(_03742_),
    .ZN(_00540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08676_ (.A1(\u_cpu.rf_ram.memory[39][6] ),
    .A2(_03738_),
    .ZN(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08677_ (.A1(_03682_),
    .A2(_03735_),
    .B(_03743_),
    .ZN(_00541_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08678_ (.A1(\u_cpu.rf_ram.memory[39][7] ),
    .A2(_03733_),
    .ZN(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08679_ (.A1(_03684_),
    .A2(_03735_),
    .B(_03744_),
    .ZN(_00542_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08680_ (.I(_03484_),
    .Z(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08681_ (.A1(_03019_),
    .A2(_03698_),
    .ZN(_03746_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08682_ (.I(_03746_),
    .Z(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08683_ (.I(_03746_),
    .Z(_03748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08684_ (.A1(\u_cpu.rf_ram.memory[137][0] ),
    .A2(_03748_),
    .ZN(_03749_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08685_ (.A1(_03745_),
    .A2(_03747_),
    .B(_03749_),
    .ZN(_00543_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08686_ (.I(_03490_),
    .Z(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08687_ (.A1(\u_cpu.rf_ram.memory[137][1] ),
    .A2(_03748_),
    .ZN(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08688_ (.A1(_03750_),
    .A2(_03747_),
    .B(_03751_),
    .ZN(_00544_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08689_ (.I(_03493_),
    .Z(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08690_ (.I(_03746_),
    .Z(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08691_ (.A1(\u_cpu.rf_ram.memory[137][2] ),
    .A2(_03753_),
    .ZN(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08692_ (.A1(_03752_),
    .A2(_03747_),
    .B(_03754_),
    .ZN(_00545_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08693_ (.I(_03497_),
    .Z(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08694_ (.A1(\u_cpu.rf_ram.memory[137][3] ),
    .A2(_03753_),
    .ZN(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08695_ (.A1(_03755_),
    .A2(_03747_),
    .B(_03756_),
    .ZN(_00546_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08696_ (.I(_03500_),
    .Z(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08697_ (.A1(\u_cpu.rf_ram.memory[137][4] ),
    .A2(_03753_),
    .ZN(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08698_ (.A1(_03757_),
    .A2(_03747_),
    .B(_03758_),
    .ZN(_00547_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08699_ (.I(_03503_),
    .Z(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08700_ (.A1(\u_cpu.rf_ram.memory[137][5] ),
    .A2(_03753_),
    .ZN(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08701_ (.A1(_03759_),
    .A2(_03748_),
    .B(_03760_),
    .ZN(_00548_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08702_ (.I(_03506_),
    .Z(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08703_ (.A1(\u_cpu.rf_ram.memory[137][6] ),
    .A2(_03753_),
    .ZN(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08704_ (.A1(_03761_),
    .A2(_03748_),
    .B(_03762_),
    .ZN(_00549_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08705_ (.I(_03509_),
    .Z(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08706_ (.A1(\u_cpu.rf_ram.memory[137][7] ),
    .A2(_03746_),
    .ZN(_03764_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08707_ (.A1(_03763_),
    .A2(_03748_),
    .B(_03764_),
    .ZN(_00550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08708_ (.A1(_02803_),
    .A2(_03380_),
    .ZN(_03765_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08709_ (.I(_03765_),
    .Z(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08710_ (.I(_03765_),
    .Z(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08711_ (.A1(\u_cpu.rf_ram.memory[49][0] ),
    .A2(_03767_),
    .ZN(_03768_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08712_ (.A1(_03745_),
    .A2(_03766_),
    .B(_03768_),
    .ZN(_00551_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08713_ (.A1(\u_cpu.rf_ram.memory[49][1] ),
    .A2(_03767_),
    .ZN(_03769_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08714_ (.A1(_03750_),
    .A2(_03766_),
    .B(_03769_),
    .ZN(_00552_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08715_ (.I(_03765_),
    .Z(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08716_ (.A1(\u_cpu.rf_ram.memory[49][2] ),
    .A2(_03770_),
    .ZN(_03771_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08717_ (.A1(_03752_),
    .A2(_03766_),
    .B(_03771_),
    .ZN(_00553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08718_ (.A1(\u_cpu.rf_ram.memory[49][3] ),
    .A2(_03770_),
    .ZN(_03772_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08719_ (.A1(_03755_),
    .A2(_03766_),
    .B(_03772_),
    .ZN(_00554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08720_ (.A1(\u_cpu.rf_ram.memory[49][4] ),
    .A2(_03770_),
    .ZN(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08721_ (.A1(_03757_),
    .A2(_03766_),
    .B(_03773_),
    .ZN(_00555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08722_ (.A1(\u_cpu.rf_ram.memory[49][5] ),
    .A2(_03770_),
    .ZN(_03774_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08723_ (.A1(_03759_),
    .A2(_03767_),
    .B(_03774_),
    .ZN(_00556_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08724_ (.A1(\u_cpu.rf_ram.memory[49][6] ),
    .A2(_03770_),
    .ZN(_03775_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08725_ (.A1(_03761_),
    .A2(_03767_),
    .B(_03775_),
    .ZN(_00557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08726_ (.A1(\u_cpu.rf_ram.memory[49][7] ),
    .A2(_03765_),
    .ZN(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08727_ (.A1(_03763_),
    .A2(_03767_),
    .B(_03776_),
    .ZN(_00558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08728_ (.A1(_03165_),
    .A2(_03698_),
    .ZN(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08729_ (.I(_03777_),
    .Z(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08730_ (.I(_03777_),
    .Z(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08731_ (.A1(\u_cpu.rf_ram.memory[136][0] ),
    .A2(_03779_),
    .ZN(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08732_ (.A1(_03745_),
    .A2(_03778_),
    .B(_03780_),
    .ZN(_00559_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08733_ (.A1(\u_cpu.rf_ram.memory[136][1] ),
    .A2(_03779_),
    .ZN(_03781_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08734_ (.A1(_03750_),
    .A2(_03778_),
    .B(_03781_),
    .ZN(_00560_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08735_ (.I(_03777_),
    .Z(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08736_ (.A1(\u_cpu.rf_ram.memory[136][2] ),
    .A2(_03782_),
    .ZN(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08737_ (.A1(_03752_),
    .A2(_03778_),
    .B(_03783_),
    .ZN(_00561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08738_ (.A1(\u_cpu.rf_ram.memory[136][3] ),
    .A2(_03782_),
    .ZN(_03784_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08739_ (.A1(_03755_),
    .A2(_03778_),
    .B(_03784_),
    .ZN(_00562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08740_ (.A1(\u_cpu.rf_ram.memory[136][4] ),
    .A2(_03782_),
    .ZN(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08741_ (.A1(_03757_),
    .A2(_03778_),
    .B(_03785_),
    .ZN(_00563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08742_ (.A1(\u_cpu.rf_ram.memory[136][5] ),
    .A2(_03782_),
    .ZN(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08743_ (.A1(_03759_),
    .A2(_03779_),
    .B(_03786_),
    .ZN(_00564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08744_ (.A1(\u_cpu.rf_ram.memory[136][6] ),
    .A2(_03782_),
    .ZN(_03787_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08745_ (.A1(_03761_),
    .A2(_03779_),
    .B(_03787_),
    .ZN(_00565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08746_ (.A1(\u_cpu.rf_ram.memory[136][7] ),
    .A2(_03777_),
    .ZN(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08747_ (.A1(_03763_),
    .A2(_03779_),
    .B(_03788_),
    .ZN(_00566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08748_ (.A1(_02876_),
    .A2(_03698_),
    .ZN(_03789_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08749_ (.I(_03789_),
    .Z(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08750_ (.I(_03789_),
    .Z(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08751_ (.A1(\u_cpu.rf_ram.memory[135][0] ),
    .A2(_03791_),
    .ZN(_03792_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08752_ (.A1(_03745_),
    .A2(_03790_),
    .B(_03792_),
    .ZN(_00567_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08753_ (.A1(\u_cpu.rf_ram.memory[135][1] ),
    .A2(_03791_),
    .ZN(_03793_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08754_ (.A1(_03750_),
    .A2(_03790_),
    .B(_03793_),
    .ZN(_00568_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08755_ (.I(_03789_),
    .Z(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08756_ (.A1(\u_cpu.rf_ram.memory[135][2] ),
    .A2(_03794_),
    .ZN(_03795_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08757_ (.A1(_03752_),
    .A2(_03790_),
    .B(_03795_),
    .ZN(_00569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08758_ (.A1(\u_cpu.rf_ram.memory[135][3] ),
    .A2(_03794_),
    .ZN(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08759_ (.A1(_03755_),
    .A2(_03790_),
    .B(_03796_),
    .ZN(_00570_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08760_ (.A1(\u_cpu.rf_ram.memory[135][4] ),
    .A2(_03794_),
    .ZN(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08761_ (.A1(_03757_),
    .A2(_03790_),
    .B(_03797_),
    .ZN(_00571_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08762_ (.A1(\u_cpu.rf_ram.memory[135][5] ),
    .A2(_03794_),
    .ZN(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08763_ (.A1(_03759_),
    .A2(_03791_),
    .B(_03798_),
    .ZN(_00572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08764_ (.A1(\u_cpu.rf_ram.memory[135][6] ),
    .A2(_03794_),
    .ZN(_03799_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08765_ (.A1(_03761_),
    .A2(_03791_),
    .B(_03799_),
    .ZN(_00573_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08766_ (.A1(\u_cpu.rf_ram.memory[135][7] ),
    .A2(_03789_),
    .ZN(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08767_ (.A1(_03763_),
    .A2(_03791_),
    .B(_03800_),
    .ZN(_00574_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08768_ (.A1(_03201_),
    .A2(_03287_),
    .ZN(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08769_ (.I(_03801_),
    .Z(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08770_ (.I(_03801_),
    .Z(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08771_ (.A1(\u_cpu.rf_ram.memory[134][0] ),
    .A2(_03803_),
    .ZN(_03804_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08772_ (.A1(_03745_),
    .A2(_03802_),
    .B(_03804_),
    .ZN(_00575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08773_ (.A1(\u_cpu.rf_ram.memory[134][1] ),
    .A2(_03803_),
    .ZN(_03805_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08774_ (.A1(_03750_),
    .A2(_03802_),
    .B(_03805_),
    .ZN(_00576_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08775_ (.I(_03801_),
    .Z(_03806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08776_ (.A1(\u_cpu.rf_ram.memory[134][2] ),
    .A2(_03806_),
    .ZN(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08777_ (.A1(_03752_),
    .A2(_03802_),
    .B(_03807_),
    .ZN(_00577_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08778_ (.A1(\u_cpu.rf_ram.memory[134][3] ),
    .A2(_03806_),
    .ZN(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08779_ (.A1(_03755_),
    .A2(_03802_),
    .B(_03808_),
    .ZN(_00578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08780_ (.A1(\u_cpu.rf_ram.memory[134][4] ),
    .A2(_03806_),
    .ZN(_03809_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08781_ (.A1(_03757_),
    .A2(_03802_),
    .B(_03809_),
    .ZN(_00579_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08782_ (.A1(\u_cpu.rf_ram.memory[134][5] ),
    .A2(_03806_),
    .ZN(_03810_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08783_ (.A1(_03759_),
    .A2(_03803_),
    .B(_03810_),
    .ZN(_00580_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08784_ (.A1(\u_cpu.rf_ram.memory[134][6] ),
    .A2(_03806_),
    .ZN(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08785_ (.A1(_03761_),
    .A2(_03803_),
    .B(_03811_),
    .ZN(_00581_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08786_ (.A1(\u_cpu.rf_ram.memory[134][7] ),
    .A2(_03801_),
    .ZN(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08787_ (.A1(_03763_),
    .A2(_03803_),
    .B(_03812_),
    .ZN(_00582_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08788_ (.I(_03484_),
    .Z(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08789_ (.I(_03201_),
    .Z(_03814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08790_ (.A1(_02786_),
    .A2(_03814_),
    .ZN(_03815_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08791_ (.I(_03815_),
    .Z(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08792_ (.I(_03815_),
    .Z(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08793_ (.A1(\u_cpu.rf_ram.memory[133][0] ),
    .A2(_03817_),
    .ZN(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08794_ (.A1(_03813_),
    .A2(_03816_),
    .B(_03818_),
    .ZN(_00583_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08795_ (.I(_03490_),
    .Z(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08796_ (.A1(\u_cpu.rf_ram.memory[133][1] ),
    .A2(_03817_),
    .ZN(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08797_ (.A1(_03819_),
    .A2(_03816_),
    .B(_03820_),
    .ZN(_00584_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08798_ (.I(_03493_),
    .Z(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08799_ (.I(_03815_),
    .Z(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08800_ (.A1(\u_cpu.rf_ram.memory[133][2] ),
    .A2(_03822_),
    .ZN(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08801_ (.A1(_03821_),
    .A2(_03816_),
    .B(_03823_),
    .ZN(_00585_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08802_ (.I(_03497_),
    .Z(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08803_ (.A1(\u_cpu.rf_ram.memory[133][3] ),
    .A2(_03822_),
    .ZN(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08804_ (.A1(_03824_),
    .A2(_03816_),
    .B(_03825_),
    .ZN(_00586_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08805_ (.I(_03500_),
    .Z(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08806_ (.A1(\u_cpu.rf_ram.memory[133][4] ),
    .A2(_03822_),
    .ZN(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08807_ (.A1(_03826_),
    .A2(_03816_),
    .B(_03827_),
    .ZN(_00587_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08808_ (.I(_03503_),
    .Z(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08809_ (.A1(\u_cpu.rf_ram.memory[133][5] ),
    .A2(_03822_),
    .ZN(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08810_ (.A1(_03828_),
    .A2(_03817_),
    .B(_03829_),
    .ZN(_00588_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08811_ (.I(_03506_),
    .Z(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08812_ (.A1(\u_cpu.rf_ram.memory[133][6] ),
    .A2(_03822_),
    .ZN(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08813_ (.A1(_03830_),
    .A2(_03817_),
    .B(_03831_),
    .ZN(_00589_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08814_ (.I(_03509_),
    .Z(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08815_ (.A1(\u_cpu.rf_ram.memory[133][7] ),
    .A2(_03815_),
    .ZN(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08816_ (.A1(_03832_),
    .A2(_03817_),
    .B(_03833_),
    .ZN(_00590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08817_ (.A1(_02830_),
    .A2(_03814_),
    .ZN(_03834_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08818_ (.I(_03834_),
    .Z(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08819_ (.I(_03834_),
    .Z(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08820_ (.A1(\u_cpu.rf_ram.memory[132][0] ),
    .A2(_03836_),
    .ZN(_03837_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08821_ (.A1(_03813_),
    .A2(_03835_),
    .B(_03837_),
    .ZN(_00591_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08822_ (.A1(\u_cpu.rf_ram.memory[132][1] ),
    .A2(_03836_),
    .ZN(_03838_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08823_ (.A1(_03819_),
    .A2(_03835_),
    .B(_03838_),
    .ZN(_00592_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08824_ (.I(_03834_),
    .Z(_03839_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08825_ (.A1(\u_cpu.rf_ram.memory[132][2] ),
    .A2(_03839_),
    .ZN(_03840_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08826_ (.A1(_03821_),
    .A2(_03835_),
    .B(_03840_),
    .ZN(_00593_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08827_ (.A1(\u_cpu.rf_ram.memory[132][3] ),
    .A2(_03839_),
    .ZN(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08828_ (.A1(_03824_),
    .A2(_03835_),
    .B(_03841_),
    .ZN(_00594_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08829_ (.A1(\u_cpu.rf_ram.memory[132][4] ),
    .A2(_03839_),
    .ZN(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08830_ (.A1(_03826_),
    .A2(_03835_),
    .B(_03842_),
    .ZN(_00595_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08831_ (.A1(\u_cpu.rf_ram.memory[132][5] ),
    .A2(_03839_),
    .ZN(_03843_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08832_ (.A1(_03828_),
    .A2(_03836_),
    .B(_03843_),
    .ZN(_00596_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08833_ (.A1(\u_cpu.rf_ram.memory[132][6] ),
    .A2(_03839_),
    .ZN(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08834_ (.A1(_03830_),
    .A2(_03836_),
    .B(_03844_),
    .ZN(_00597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08835_ (.A1(\u_cpu.rf_ram.memory[132][7] ),
    .A2(_03834_),
    .ZN(_03845_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08836_ (.A1(_03832_),
    .A2(_03836_),
    .B(_03845_),
    .ZN(_00598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08837_ (.A1(_03002_),
    .A2(_03814_),
    .ZN(_03846_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08838_ (.I(_03846_),
    .Z(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08839_ (.I(_03846_),
    .Z(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08840_ (.A1(\u_cpu.rf_ram.memory[131][0] ),
    .A2(_03848_),
    .ZN(_03849_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08841_ (.A1(_03813_),
    .A2(_03847_),
    .B(_03849_),
    .ZN(_00599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08842_ (.A1(\u_cpu.rf_ram.memory[131][1] ),
    .A2(_03848_),
    .ZN(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08843_ (.A1(_03819_),
    .A2(_03847_),
    .B(_03850_),
    .ZN(_00600_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08844_ (.I(_03846_),
    .Z(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08845_ (.A1(\u_cpu.rf_ram.memory[131][2] ),
    .A2(_03851_),
    .ZN(_03852_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08846_ (.A1(_03821_),
    .A2(_03847_),
    .B(_03852_),
    .ZN(_00601_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08847_ (.A1(\u_cpu.rf_ram.memory[131][3] ),
    .A2(_03851_),
    .ZN(_03853_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08848_ (.A1(_03824_),
    .A2(_03847_),
    .B(_03853_),
    .ZN(_00602_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08849_ (.A1(\u_cpu.rf_ram.memory[131][4] ),
    .A2(_03851_),
    .ZN(_03854_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08850_ (.A1(_03826_),
    .A2(_03847_),
    .B(_03854_),
    .ZN(_00603_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08851_ (.A1(\u_cpu.rf_ram.memory[131][5] ),
    .A2(_03851_),
    .ZN(_03855_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08852_ (.A1(_03828_),
    .A2(_03848_),
    .B(_03855_),
    .ZN(_00604_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08853_ (.A1(\u_cpu.rf_ram.memory[131][6] ),
    .A2(_03851_),
    .ZN(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08854_ (.A1(_03830_),
    .A2(_03848_),
    .B(_03856_),
    .ZN(_00605_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08855_ (.A1(\u_cpu.rf_ram.memory[131][7] ),
    .A2(_03846_),
    .ZN(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08856_ (.A1(_03832_),
    .A2(_03848_),
    .B(_03857_),
    .ZN(_00606_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08857_ (.A1(_02722_),
    .A2(_03814_),
    .ZN(_03858_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08858_ (.I(_03858_),
    .Z(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08859_ (.I(_03858_),
    .Z(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08860_ (.A1(\u_cpu.rf_ram.memory[130][0] ),
    .A2(_03860_),
    .ZN(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08861_ (.A1(_03813_),
    .A2(_03859_),
    .B(_03861_),
    .ZN(_00607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08862_ (.A1(\u_cpu.rf_ram.memory[130][1] ),
    .A2(_03860_),
    .ZN(_03862_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08863_ (.A1(_03819_),
    .A2(_03859_),
    .B(_03862_),
    .ZN(_00608_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08864_ (.I(_03858_),
    .Z(_03863_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08865_ (.A1(\u_cpu.rf_ram.memory[130][2] ),
    .A2(_03863_),
    .ZN(_03864_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08866_ (.A1(_03821_),
    .A2(_03859_),
    .B(_03864_),
    .ZN(_00609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08867_ (.A1(\u_cpu.rf_ram.memory[130][3] ),
    .A2(_03863_),
    .ZN(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08868_ (.A1(_03824_),
    .A2(_03859_),
    .B(_03865_),
    .ZN(_00610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08869_ (.A1(\u_cpu.rf_ram.memory[130][4] ),
    .A2(_03863_),
    .ZN(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08870_ (.A1(_03826_),
    .A2(_03859_),
    .B(_03866_),
    .ZN(_00611_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08871_ (.A1(\u_cpu.rf_ram.memory[130][5] ),
    .A2(_03863_),
    .ZN(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08872_ (.A1(_03828_),
    .A2(_03860_),
    .B(_03867_),
    .ZN(_00612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08873_ (.A1(\u_cpu.rf_ram.memory[130][6] ),
    .A2(_03863_),
    .ZN(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08874_ (.A1(_03830_),
    .A2(_03860_),
    .B(_03868_),
    .ZN(_00613_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08875_ (.A1(\u_cpu.rf_ram.memory[130][7] ),
    .A2(_03858_),
    .ZN(_03869_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08876_ (.A1(_03832_),
    .A2(_03860_),
    .B(_03869_),
    .ZN(_00614_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08877_ (.I(_02849_),
    .Z(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08878_ (.A1(_03870_),
    .A2(_02982_),
    .ZN(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08879_ (.I(_03871_),
    .Z(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08880_ (.I0(_03560_),
    .I1(\u_cpu.rf_ram.memory[12][0] ),
    .S(_03872_),
    .Z(_03873_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08881_ (.I(_03873_),
    .Z(_00615_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08882_ (.I0(_03564_),
    .I1(\u_cpu.rf_ram.memory[12][1] ),
    .S(_03872_),
    .Z(_03874_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08883_ (.I(_03874_),
    .Z(_00616_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08884_ (.I0(_03566_),
    .I1(\u_cpu.rf_ram.memory[12][2] ),
    .S(_03872_),
    .Z(_03875_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08885_ (.I(_03875_),
    .Z(_00617_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08886_ (.I0(_03568_),
    .I1(\u_cpu.rf_ram.memory[12][3] ),
    .S(_03872_),
    .Z(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08887_ (.I(_03876_),
    .Z(_00618_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08888_ (.I0(_03570_),
    .I1(\u_cpu.rf_ram.memory[12][4] ),
    .S(_03872_),
    .Z(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08889_ (.I(_03877_),
    .Z(_00619_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08890_ (.I0(_03572_),
    .I1(\u_cpu.rf_ram.memory[12][5] ),
    .S(_03871_),
    .Z(_03878_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08891_ (.I(_03878_),
    .Z(_00620_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08892_ (.I0(_03574_),
    .I1(\u_cpu.rf_ram.memory[12][6] ),
    .S(_03871_),
    .Z(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08893_ (.I(_03879_),
    .Z(_00621_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08894_ (.I0(_03576_),
    .I1(\u_cpu.rf_ram.memory[12][7] ),
    .S(_03871_),
    .Z(_03880_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08895_ (.I(_03880_),
    .Z(_00622_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08896_ (.A1(_03367_),
    .A2(_03287_),
    .ZN(_03881_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08897_ (.I(_03881_),
    .Z(_03882_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08898_ (.I(_03881_),
    .Z(_03883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08899_ (.A1(\u_cpu.rf_ram.memory[22][0] ),
    .A2(_03883_),
    .ZN(_03884_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08900_ (.A1(_03813_),
    .A2(_03882_),
    .B(_03884_),
    .ZN(_00623_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08901_ (.A1(\u_cpu.rf_ram.memory[22][1] ),
    .A2(_03883_),
    .ZN(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08902_ (.A1(_03819_),
    .A2(_03882_),
    .B(_03885_),
    .ZN(_00624_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08903_ (.I(_03881_),
    .Z(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08904_ (.A1(\u_cpu.rf_ram.memory[22][2] ),
    .A2(_03886_),
    .ZN(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08905_ (.A1(_03821_),
    .A2(_03882_),
    .B(_03887_),
    .ZN(_00625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08906_ (.A1(\u_cpu.rf_ram.memory[22][3] ),
    .A2(_03886_),
    .ZN(_03888_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08907_ (.A1(_03824_),
    .A2(_03882_),
    .B(_03888_),
    .ZN(_00626_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08908_ (.A1(\u_cpu.rf_ram.memory[22][4] ),
    .A2(_03886_),
    .ZN(_03889_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08909_ (.A1(_03826_),
    .A2(_03882_),
    .B(_03889_),
    .ZN(_00627_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08910_ (.A1(\u_cpu.rf_ram.memory[22][5] ),
    .A2(_03886_),
    .ZN(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08911_ (.A1(_03828_),
    .A2(_03883_),
    .B(_03890_),
    .ZN(_00628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08912_ (.A1(\u_cpu.rf_ram.memory[22][6] ),
    .A2(_03886_),
    .ZN(_03891_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08913_ (.A1(_03830_),
    .A2(_03883_),
    .B(_03891_),
    .ZN(_00629_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08914_ (.A1(\u_cpu.rf_ram.memory[22][7] ),
    .A2(_03881_),
    .ZN(_03892_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08915_ (.A1(_03832_),
    .A2(_03883_),
    .B(_03892_),
    .ZN(_00630_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08916_ (.I(_02738_),
    .Z(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08917_ (.I(_03893_),
    .Z(_03894_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08918_ (.A1(_02890_),
    .A2(_03814_),
    .ZN(_03895_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08919_ (.I(_03895_),
    .Z(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08920_ (.I(_03895_),
    .Z(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08921_ (.A1(\u_cpu.rf_ram.memory[128][0] ),
    .A2(_03897_),
    .ZN(_03898_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08922_ (.A1(_03894_),
    .A2(_03896_),
    .B(_03898_),
    .ZN(_00631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08923_ (.I(_02744_),
    .Z(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08924_ (.I(_03899_),
    .Z(_03900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08925_ (.A1(\u_cpu.rf_ram.memory[128][1] ),
    .A2(_03897_),
    .ZN(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08926_ (.A1(_03900_),
    .A2(_03896_),
    .B(_03901_),
    .ZN(_00632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08927_ (.I(_02750_),
    .Z(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08928_ (.I(_03902_),
    .Z(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08929_ (.I(_03895_),
    .Z(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08930_ (.A1(\u_cpu.rf_ram.memory[128][2] ),
    .A2(_03904_),
    .ZN(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08931_ (.A1(_03903_),
    .A2(_03896_),
    .B(_03905_),
    .ZN(_00633_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08932_ (.I(_02756_),
    .Z(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08933_ (.I(_03906_),
    .Z(_03907_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08934_ (.A1(\u_cpu.rf_ram.memory[128][3] ),
    .A2(_03904_),
    .ZN(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08935_ (.A1(_03907_),
    .A2(_03896_),
    .B(_03908_),
    .ZN(_00634_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08936_ (.I(_02761_),
    .Z(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08937_ (.I(_03909_),
    .Z(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08938_ (.A1(\u_cpu.rf_ram.memory[128][4] ),
    .A2(_03904_),
    .ZN(_03911_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08939_ (.A1(_03910_),
    .A2(_03896_),
    .B(_03911_),
    .ZN(_00635_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08940_ (.I(_02766_),
    .Z(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08941_ (.I(_03912_),
    .Z(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08942_ (.A1(\u_cpu.rf_ram.memory[128][5] ),
    .A2(_03904_),
    .ZN(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08943_ (.A1(_03913_),
    .A2(_03897_),
    .B(_03914_),
    .ZN(_00636_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08944_ (.I(_02771_),
    .Z(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08945_ (.I(_03915_),
    .Z(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08946_ (.A1(\u_cpu.rf_ram.memory[128][6] ),
    .A2(_03904_),
    .ZN(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08947_ (.A1(_03916_),
    .A2(_03897_),
    .B(_03917_),
    .ZN(_00637_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08948_ (.I(_02776_),
    .Z(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08949_ (.I(_03918_),
    .Z(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08950_ (.A1(\u_cpu.rf_ram.memory[128][7] ),
    .A2(_03895_),
    .ZN(_03920_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08951_ (.A1(_03919_),
    .A2(_03897_),
    .B(_03920_),
    .ZN(_00638_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08952_ (.A1(_03061_),
    .A2(_03181_),
    .ZN(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08953_ (.I(_03921_),
    .Z(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08954_ (.I(_03921_),
    .Z(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08955_ (.A1(\u_cpu.rf_ram.memory[127][0] ),
    .A2(_03923_),
    .ZN(_03924_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08956_ (.A1(_03894_),
    .A2(_03922_),
    .B(_03924_),
    .ZN(_00639_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08957_ (.A1(\u_cpu.rf_ram.memory[127][1] ),
    .A2(_03923_),
    .ZN(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08958_ (.A1(_03900_),
    .A2(_03922_),
    .B(_03925_),
    .ZN(_00640_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08959_ (.I(_03921_),
    .Z(_03926_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08960_ (.A1(\u_cpu.rf_ram.memory[127][2] ),
    .A2(_03926_),
    .ZN(_03927_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08961_ (.A1(_03903_),
    .A2(_03922_),
    .B(_03927_),
    .ZN(_00641_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08962_ (.A1(\u_cpu.rf_ram.memory[127][3] ),
    .A2(_03926_),
    .ZN(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08963_ (.A1(_03907_),
    .A2(_03922_),
    .B(_03928_),
    .ZN(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08964_ (.A1(\u_cpu.rf_ram.memory[127][4] ),
    .A2(_03926_),
    .ZN(_03929_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08965_ (.A1(_03910_),
    .A2(_03922_),
    .B(_03929_),
    .ZN(_00643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08966_ (.A1(\u_cpu.rf_ram.memory[127][5] ),
    .A2(_03926_),
    .ZN(_03930_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08967_ (.A1(_03913_),
    .A2(_03923_),
    .B(_03930_),
    .ZN(_00644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08968_ (.A1(\u_cpu.rf_ram.memory[127][6] ),
    .A2(_03926_),
    .ZN(_03931_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08969_ (.A1(_03916_),
    .A2(_03923_),
    .B(_03931_),
    .ZN(_00645_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08970_ (.A1(\u_cpu.rf_ram.memory[127][7] ),
    .A2(_03921_),
    .ZN(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08971_ (.A1(_03919_),
    .A2(_03923_),
    .B(_03932_),
    .ZN(_00646_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08972_ (.A1(_02920_),
    .A2(_03181_),
    .ZN(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08973_ (.I(_03933_),
    .Z(_03934_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08974_ (.I(_03933_),
    .Z(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08975_ (.A1(\u_cpu.rf_ram.memory[126][0] ),
    .A2(_03935_),
    .ZN(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08976_ (.A1(_03894_),
    .A2(_03934_),
    .B(_03936_),
    .ZN(_00647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08977_ (.A1(\u_cpu.rf_ram.memory[126][1] ),
    .A2(_03935_),
    .ZN(_03937_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08978_ (.A1(_03900_),
    .A2(_03934_),
    .B(_03937_),
    .ZN(_00648_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08979_ (.I(_03933_),
    .Z(_03938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08980_ (.A1(\u_cpu.rf_ram.memory[126][2] ),
    .A2(_03938_),
    .ZN(_03939_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08981_ (.A1(_03903_),
    .A2(_03934_),
    .B(_03939_),
    .ZN(_00649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08982_ (.A1(\u_cpu.rf_ram.memory[126][3] ),
    .A2(_03938_),
    .ZN(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08983_ (.A1(_03907_),
    .A2(_03934_),
    .B(_03940_),
    .ZN(_00650_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08984_ (.A1(\u_cpu.rf_ram.memory[126][4] ),
    .A2(_03938_),
    .ZN(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08985_ (.A1(_03910_),
    .A2(_03934_),
    .B(_03941_),
    .ZN(_00651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08986_ (.A1(\u_cpu.rf_ram.memory[126][5] ),
    .A2(_03938_),
    .ZN(_03942_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08987_ (.A1(_03913_),
    .A2(_03935_),
    .B(_03942_),
    .ZN(_00652_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08988_ (.A1(\u_cpu.rf_ram.memory[126][6] ),
    .A2(_03938_),
    .ZN(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08989_ (.A1(_03916_),
    .A2(_03935_),
    .B(_03943_),
    .ZN(_00653_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08990_ (.A1(\u_cpu.rf_ram.memory[126][7] ),
    .A2(_03933_),
    .ZN(_03944_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08991_ (.A1(_03919_),
    .A2(_03935_),
    .B(_03944_),
    .ZN(_00654_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08992_ (.A1(_02966_),
    .A2(_03181_),
    .ZN(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08993_ (.I(_03945_),
    .Z(_03946_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08994_ (.I(_03945_),
    .Z(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08995_ (.A1(\u_cpu.rf_ram.memory[125][0] ),
    .A2(_03947_),
    .ZN(_03948_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08996_ (.A1(_03894_),
    .A2(_03946_),
    .B(_03948_),
    .ZN(_00655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08997_ (.A1(\u_cpu.rf_ram.memory[125][1] ),
    .A2(_03947_),
    .ZN(_03949_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08998_ (.A1(_03900_),
    .A2(_03946_),
    .B(_03949_),
    .ZN(_00656_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08999_ (.I(_03945_),
    .Z(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09000_ (.A1(\u_cpu.rf_ram.memory[125][2] ),
    .A2(_03950_),
    .ZN(_03951_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09001_ (.A1(_03903_),
    .A2(_03946_),
    .B(_03951_),
    .ZN(_00657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09002_ (.A1(\u_cpu.rf_ram.memory[125][3] ),
    .A2(_03950_),
    .ZN(_03952_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09003_ (.A1(_03907_),
    .A2(_03946_),
    .B(_03952_),
    .ZN(_00658_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09004_ (.A1(\u_cpu.rf_ram.memory[125][4] ),
    .A2(_03950_),
    .ZN(_03953_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09005_ (.A1(_03910_),
    .A2(_03946_),
    .B(_03953_),
    .ZN(_00659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09006_ (.A1(\u_cpu.rf_ram.memory[125][5] ),
    .A2(_03950_),
    .ZN(_03954_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09007_ (.A1(_03913_),
    .A2(_03947_),
    .B(_03954_),
    .ZN(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09008_ (.A1(\u_cpu.rf_ram.memory[125][6] ),
    .A2(_03950_),
    .ZN(_03955_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09009_ (.A1(_03916_),
    .A2(_03947_),
    .B(_03955_),
    .ZN(_00661_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09010_ (.A1(\u_cpu.rf_ram.memory[125][7] ),
    .A2(_03945_),
    .ZN(_03956_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09011_ (.A1(_03919_),
    .A2(_03947_),
    .B(_03956_),
    .ZN(_00662_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09012_ (.A1(_02981_),
    .A2(_03181_),
    .ZN(_03957_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09013_ (.I(_03957_),
    .Z(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09014_ (.I(_03957_),
    .Z(_03959_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09015_ (.A1(\u_cpu.rf_ram.memory[124][0] ),
    .A2(_03959_),
    .ZN(_03960_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09016_ (.A1(_03894_),
    .A2(_03958_),
    .B(_03960_),
    .ZN(_00663_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09017_ (.A1(\u_cpu.rf_ram.memory[124][1] ),
    .A2(_03959_),
    .ZN(_03961_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09018_ (.A1(_03900_),
    .A2(_03958_),
    .B(_03961_),
    .ZN(_00664_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09019_ (.I(_03957_),
    .Z(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09020_ (.A1(\u_cpu.rf_ram.memory[124][2] ),
    .A2(_03962_),
    .ZN(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09021_ (.A1(_03903_),
    .A2(_03958_),
    .B(_03963_),
    .ZN(_00665_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09022_ (.A1(\u_cpu.rf_ram.memory[124][3] ),
    .A2(_03962_),
    .ZN(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09023_ (.A1(_03907_),
    .A2(_03958_),
    .B(_03964_),
    .ZN(_00666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09024_ (.A1(\u_cpu.rf_ram.memory[124][4] ),
    .A2(_03962_),
    .ZN(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09025_ (.A1(_03910_),
    .A2(_03958_),
    .B(_03965_),
    .ZN(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09026_ (.A1(\u_cpu.rf_ram.memory[124][5] ),
    .A2(_03962_),
    .ZN(_03966_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09027_ (.A1(_03913_),
    .A2(_03959_),
    .B(_03966_),
    .ZN(_00668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09028_ (.A1(\u_cpu.rf_ram.memory[124][6] ),
    .A2(_03962_),
    .ZN(_03967_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09029_ (.A1(_03916_),
    .A2(_03959_),
    .B(_03967_),
    .ZN(_00669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09030_ (.A1(\u_cpu.rf_ram.memory[124][7] ),
    .A2(_03957_),
    .ZN(_03968_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09031_ (.A1(_03919_),
    .A2(_03959_),
    .B(_03968_),
    .ZN(_00670_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09032_ (.I(_03893_),
    .Z(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09033_ (.I(_03180_),
    .Z(_03970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09034_ (.A1(_03033_),
    .A2(_03970_),
    .ZN(_03971_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09035_ (.I(_03971_),
    .Z(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09036_ (.I(_03971_),
    .Z(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09037_ (.A1(\u_cpu.rf_ram.memory[123][0] ),
    .A2(_03973_),
    .ZN(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09038_ (.A1(_03969_),
    .A2(_03972_),
    .B(_03974_),
    .ZN(_00671_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09039_ (.I(_03899_),
    .Z(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09040_ (.A1(\u_cpu.rf_ram.memory[123][1] ),
    .A2(_03973_),
    .ZN(_03976_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09041_ (.A1(_03975_),
    .A2(_03972_),
    .B(_03976_),
    .ZN(_00672_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09042_ (.I(_03902_),
    .Z(_03977_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09043_ (.I(_03971_),
    .Z(_03978_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09044_ (.A1(\u_cpu.rf_ram.memory[123][2] ),
    .A2(_03978_),
    .ZN(_03979_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09045_ (.A1(_03977_),
    .A2(_03972_),
    .B(_03979_),
    .ZN(_00673_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09046_ (.I(_03906_),
    .Z(_03980_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09047_ (.A1(\u_cpu.rf_ram.memory[123][3] ),
    .A2(_03978_),
    .ZN(_03981_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09048_ (.A1(_03980_),
    .A2(_03972_),
    .B(_03981_),
    .ZN(_00674_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09049_ (.I(_03909_),
    .Z(_03982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09050_ (.A1(\u_cpu.rf_ram.memory[123][4] ),
    .A2(_03978_),
    .ZN(_03983_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09051_ (.A1(_03982_),
    .A2(_03972_),
    .B(_03983_),
    .ZN(_00675_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09052_ (.I(_03912_),
    .Z(_03984_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09053_ (.A1(\u_cpu.rf_ram.memory[123][5] ),
    .A2(_03978_),
    .ZN(_03985_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09054_ (.A1(_03984_),
    .A2(_03973_),
    .B(_03985_),
    .ZN(_00676_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09055_ (.I(_03915_),
    .Z(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09056_ (.A1(\u_cpu.rf_ram.memory[123][6] ),
    .A2(_03978_),
    .ZN(_03987_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09057_ (.A1(_03986_),
    .A2(_03973_),
    .B(_03987_),
    .ZN(_00677_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09058_ (.I(_03918_),
    .Z(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09059_ (.A1(\u_cpu.rf_ram.memory[123][7] ),
    .A2(_03971_),
    .ZN(_03989_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09060_ (.A1(_03988_),
    .A2(_03973_),
    .B(_03989_),
    .ZN(_00678_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09061_ (.A1(_03018_),
    .A2(_03286_),
    .ZN(_03990_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09062_ (.I(_03990_),
    .Z(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09063_ (.I(_03990_),
    .Z(_03992_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09064_ (.A1(\u_cpu.rf_ram.memory[38][0] ),
    .A2(_03992_),
    .ZN(_03993_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09065_ (.A1(_03969_),
    .A2(_03991_),
    .B(_03993_),
    .ZN(_00679_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09066_ (.A1(\u_cpu.rf_ram.memory[38][1] ),
    .A2(_03992_),
    .ZN(_03994_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09067_ (.A1(_03975_),
    .A2(_03991_),
    .B(_03994_),
    .ZN(_00680_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09068_ (.I(_03990_),
    .Z(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09069_ (.A1(\u_cpu.rf_ram.memory[38][2] ),
    .A2(_03995_),
    .ZN(_03996_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09070_ (.A1(_03977_),
    .A2(_03991_),
    .B(_03996_),
    .ZN(_00681_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09071_ (.A1(\u_cpu.rf_ram.memory[38][3] ),
    .A2(_03995_),
    .ZN(_03997_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09072_ (.A1(_03980_),
    .A2(_03991_),
    .B(_03997_),
    .ZN(_00682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09073_ (.A1(\u_cpu.rf_ram.memory[38][4] ),
    .A2(_03995_),
    .ZN(_03998_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09074_ (.A1(_03982_),
    .A2(_03991_),
    .B(_03998_),
    .ZN(_00683_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09075_ (.A1(\u_cpu.rf_ram.memory[38][5] ),
    .A2(_03995_),
    .ZN(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09076_ (.A1(_03984_),
    .A2(_03992_),
    .B(_03999_),
    .ZN(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09077_ (.A1(\u_cpu.rf_ram.memory[38][6] ),
    .A2(_03995_),
    .ZN(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09078_ (.A1(_03986_),
    .A2(_03992_),
    .B(_04000_),
    .ZN(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09079_ (.A1(\u_cpu.rf_ram.memory[38][7] ),
    .A2(_03990_),
    .ZN(_04001_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09080_ (.A1(_03988_),
    .A2(_03992_),
    .B(_04001_),
    .ZN(_00686_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09081_ (.A1(_02785_),
    .A2(_02940_),
    .ZN(_04002_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09082_ (.I(_04002_),
    .Z(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09083_ (.I(_04002_),
    .Z(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09084_ (.A1(\u_cpu.rf_ram.memory[37][0] ),
    .A2(_04004_),
    .ZN(_04005_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09085_ (.A1(_03969_),
    .A2(_04003_),
    .B(_04005_),
    .ZN(_00687_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09086_ (.A1(\u_cpu.rf_ram.memory[37][1] ),
    .A2(_04004_),
    .ZN(_04006_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09087_ (.A1(_03975_),
    .A2(_04003_),
    .B(_04006_),
    .ZN(_00688_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09088_ (.I(_04002_),
    .Z(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09089_ (.A1(\u_cpu.rf_ram.memory[37][2] ),
    .A2(_04007_),
    .ZN(_04008_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09090_ (.A1(_03977_),
    .A2(_04003_),
    .B(_04008_),
    .ZN(_00689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09091_ (.A1(\u_cpu.rf_ram.memory[37][3] ),
    .A2(_04007_),
    .ZN(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09092_ (.A1(_03980_),
    .A2(_04003_),
    .B(_04009_),
    .ZN(_00690_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09093_ (.A1(\u_cpu.rf_ram.memory[37][4] ),
    .A2(_04007_),
    .ZN(_04010_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09094_ (.A1(_03982_),
    .A2(_04003_),
    .B(_04010_),
    .ZN(_00691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09095_ (.A1(\u_cpu.rf_ram.memory[37][5] ),
    .A2(_04007_),
    .ZN(_04011_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09096_ (.A1(_03984_),
    .A2(_04004_),
    .B(_04011_),
    .ZN(_00692_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09097_ (.A1(\u_cpu.rf_ram.memory[37][6] ),
    .A2(_04007_),
    .ZN(_04012_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09098_ (.A1(_03986_),
    .A2(_04004_),
    .B(_04012_),
    .ZN(_00693_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09099_ (.A1(\u_cpu.rf_ram.memory[37][7] ),
    .A2(_04002_),
    .ZN(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09100_ (.A1(_03988_),
    .A2(_04004_),
    .B(_04013_),
    .ZN(_00694_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09101_ (.A1(_02830_),
    .A2(_02940_),
    .ZN(_04014_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09102_ (.I(_04014_),
    .Z(_04015_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09103_ (.I(_04014_),
    .Z(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09104_ (.A1(\u_cpu.rf_ram.memory[36][0] ),
    .A2(_04016_),
    .ZN(_04017_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09105_ (.A1(_03969_),
    .A2(_04015_),
    .B(_04017_),
    .ZN(_00695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09106_ (.A1(\u_cpu.rf_ram.memory[36][1] ),
    .A2(_04016_),
    .ZN(_04018_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09107_ (.A1(_03975_),
    .A2(_04015_),
    .B(_04018_),
    .ZN(_00696_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09108_ (.I(_04014_),
    .Z(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09109_ (.A1(\u_cpu.rf_ram.memory[36][2] ),
    .A2(_04019_),
    .ZN(_04020_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09110_ (.A1(_03977_),
    .A2(_04015_),
    .B(_04020_),
    .ZN(_00697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09111_ (.A1(\u_cpu.rf_ram.memory[36][3] ),
    .A2(_04019_),
    .ZN(_04021_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09112_ (.A1(_03980_),
    .A2(_04015_),
    .B(_04021_),
    .ZN(_00698_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09113_ (.A1(\u_cpu.rf_ram.memory[36][4] ),
    .A2(_04019_),
    .ZN(_04022_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09114_ (.A1(_03982_),
    .A2(_04015_),
    .B(_04022_),
    .ZN(_00699_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09115_ (.A1(\u_cpu.rf_ram.memory[36][5] ),
    .A2(_04019_),
    .ZN(_04023_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09116_ (.A1(_03984_),
    .A2(_04016_),
    .B(_04023_),
    .ZN(_00700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09117_ (.A1(\u_cpu.rf_ram.memory[36][6] ),
    .A2(_04019_),
    .ZN(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09118_ (.A1(_03986_),
    .A2(_04016_),
    .B(_04024_),
    .ZN(_00701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09119_ (.A1(\u_cpu.rf_ram.memory[36][7] ),
    .A2(_04014_),
    .ZN(_04025_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09120_ (.A1(_03988_),
    .A2(_04016_),
    .B(_04025_),
    .ZN(_00702_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09121_ (.I(_02569_),
    .Z(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09122_ (.A1(_04026_),
    .A2(_03123_),
    .ZN(_04027_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09123_ (.A1(_03111_),
    .A2(_04027_),
    .ZN(_04028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09124_ (.I(_04028_),
    .Z(_00703_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09125_ (.A1(\u_cpu.cpu.state.o_cnt[2] ),
    .A2(_02563_),
    .ZN(_04029_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09126_ (.A1(\u_cpu.cpu.state.o_cnt[2] ),
    .A2(_02563_),
    .Z(_04030_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09127_ (.A1(_03111_),
    .A2(_04029_),
    .A3(_04030_),
    .ZN(_00704_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09128_ (.I(\u_cpu.cpu.mem_bytecnt[0] ),
    .Z(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09129_ (.I(_01432_),
    .Z(_04032_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09130_ (.A1(_04031_),
    .A2(_04030_),
    .B(_04032_),
    .ZN(_04033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09131_ (.A1(_04031_),
    .A2(_04030_),
    .B(_04033_),
    .ZN(_00705_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09132_ (.I(\u_cpu.cpu.mem_bytecnt[1] ),
    .Z(_04034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09133_ (.A1(_04031_),
    .A2(_04030_),
    .ZN(_04035_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09134_ (.A1(_04034_),
    .A2(_04035_),
    .Z(_04036_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09135_ (.A1(_03112_),
    .A2(_04036_),
    .ZN(_00706_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09136_ (.A1(net2),
    .A2(_04026_),
    .ZN(_04037_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09137_ (.I(_04037_),
    .Z(_04038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09138_ (.A1(_02563_),
    .A2(_04038_),
    .ZN(_04039_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09139_ (.I(_03134_),
    .ZN(_04040_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09140_ (.A1(\u_cpu.rf_ram_if.rgnt ),
    .A2(_04040_),
    .B(_02699_),
    .C(_04032_),
    .ZN(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09141_ (.A1(_04039_),
    .A2(_04041_),
    .ZN(_00707_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09142_ (.A1(_04032_),
    .A2(\u_cpu.cpu.state.o_cnt_r[0] ),
    .Z(_04042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09143_ (.I(_04042_),
    .Z(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09144_ (.A1(_03112_),
    .A2(_02607_),
    .ZN(_00709_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09145_ (.A1(_01432_),
    .A2(\u_cpu.cpu.state.o_cnt_r[2] ),
    .Z(_04043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09146_ (.I(_04043_),
    .Z(_00710_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09147_ (.A1(_02731_),
    .A2(_03034_),
    .ZN(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09148_ (.I(_04044_),
    .Z(_04045_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09149_ (.I(_04044_),
    .Z(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09150_ (.A1(\u_cpu.rf_ram.memory[91][0] ),
    .A2(_04046_),
    .ZN(_04047_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09151_ (.A1(_03969_),
    .A2(_04045_),
    .B(_04047_),
    .ZN(_00711_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09152_ (.A1(\u_cpu.rf_ram.memory[91][1] ),
    .A2(_04046_),
    .ZN(_04048_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09153_ (.A1(_03975_),
    .A2(_04045_),
    .B(_04048_),
    .ZN(_00712_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09154_ (.I(_04044_),
    .Z(_04049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09155_ (.A1(\u_cpu.rf_ram.memory[91][2] ),
    .A2(_04049_),
    .ZN(_04050_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09156_ (.A1(_03977_),
    .A2(_04045_),
    .B(_04050_),
    .ZN(_00713_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09157_ (.A1(\u_cpu.rf_ram.memory[91][3] ),
    .A2(_04049_),
    .ZN(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09158_ (.A1(_03980_),
    .A2(_04045_),
    .B(_04051_),
    .ZN(_00714_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09159_ (.A1(\u_cpu.rf_ram.memory[91][4] ),
    .A2(_04049_),
    .ZN(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09160_ (.A1(_03982_),
    .A2(_04045_),
    .B(_04052_),
    .ZN(_00715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09161_ (.A1(\u_cpu.rf_ram.memory[91][5] ),
    .A2(_04049_),
    .ZN(_04053_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09162_ (.A1(_03984_),
    .A2(_04046_),
    .B(_04053_),
    .ZN(_00716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09163_ (.A1(\u_cpu.rf_ram.memory[91][6] ),
    .A2(_04049_),
    .ZN(_04054_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09164_ (.A1(_03986_),
    .A2(_04046_),
    .B(_04054_),
    .ZN(_00717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09165_ (.A1(\u_cpu.rf_ram.memory[91][7] ),
    .A2(_04044_),
    .ZN(_04055_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09166_ (.A1(_03988_),
    .A2(_04046_),
    .B(_04055_),
    .ZN(_00718_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09167_ (.I(_03893_),
    .Z(_04056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09168_ (.A1(_02731_),
    .A2(_02938_),
    .ZN(_04057_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09169_ (.I(_04057_),
    .Z(_04058_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09170_ (.I(_04057_),
    .Z(_04059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09171_ (.A1(\u_cpu.rf_ram.memory[90][0] ),
    .A2(_04059_),
    .ZN(_04060_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09172_ (.A1(_04056_),
    .A2(_04058_),
    .B(_04060_),
    .ZN(_00719_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09173_ (.I(_03899_),
    .Z(_04061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09174_ (.A1(\u_cpu.rf_ram.memory[90][1] ),
    .A2(_04059_),
    .ZN(_04062_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09175_ (.A1(_04061_),
    .A2(_04058_),
    .B(_04062_),
    .ZN(_00720_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09176_ (.I(_03902_),
    .Z(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09177_ (.I(_04057_),
    .Z(_04064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09178_ (.A1(\u_cpu.rf_ram.memory[90][2] ),
    .A2(_04064_),
    .ZN(_04065_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09179_ (.A1(_04063_),
    .A2(_04058_),
    .B(_04065_),
    .ZN(_00721_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09180_ (.I(_03906_),
    .Z(_04066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09181_ (.A1(\u_cpu.rf_ram.memory[90][3] ),
    .A2(_04064_),
    .ZN(_04067_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09182_ (.A1(_04066_),
    .A2(_04058_),
    .B(_04067_),
    .ZN(_00722_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09183_ (.I(_03909_),
    .Z(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09184_ (.A1(\u_cpu.rf_ram.memory[90][4] ),
    .A2(_04064_),
    .ZN(_04069_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09185_ (.A1(_04068_),
    .A2(_04058_),
    .B(_04069_),
    .ZN(_00723_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09186_ (.I(_03912_),
    .Z(_04070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09187_ (.A1(\u_cpu.rf_ram.memory[90][5] ),
    .A2(_04064_),
    .ZN(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09188_ (.A1(_04070_),
    .A2(_04059_),
    .B(_04071_),
    .ZN(_00724_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09189_ (.I(_03915_),
    .Z(_04072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09190_ (.A1(\u_cpu.rf_ram.memory[90][6] ),
    .A2(_04064_),
    .ZN(_04073_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09191_ (.A1(_04072_),
    .A2(_04059_),
    .B(_04073_),
    .ZN(_00725_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09192_ (.I(_03918_),
    .Z(_04074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09193_ (.A1(\u_cpu.rf_ram.memory[90][7] ),
    .A2(_04057_),
    .ZN(_04075_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09194_ (.A1(_04074_),
    .A2(_04059_),
    .B(_04075_),
    .ZN(_00726_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09195_ (.A1(_02673_),
    .A2(_02677_),
    .ZN(_04076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09196_ (.A1(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ),
    .A2(_04038_),
    .ZN(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09197_ (.A1(_03111_),
    .A2(_04027_),
    .A3(_04076_),
    .B(_04077_),
    .ZN(_00727_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09198_ (.A1(\u_cpu.cpu.ctrl.i_jump ),
    .A2(_04038_),
    .ZN(_04078_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09199_ (.A1(_02558_),
    .A2(_02594_),
    .ZN(_04079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09200_ (.A1(_02549_),
    .A2(_04079_),
    .ZN(_04080_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09201_ (.A1(_02547_),
    .A2(_04079_),
    .Z(_04081_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09202_ (.A1(_02551_),
    .A2(_04081_),
    .Z(_04082_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09203_ (.A1(_04080_),
    .A2(_04082_),
    .Z(_04083_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09204_ (.A1(_01409_),
    .A2(_02556_),
    .B1(_04080_),
    .B2(_04082_),
    .ZN(_04084_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09205_ (.A1(_02585_),
    .A2(_02586_),
    .B(_02553_),
    .C(_02559_),
    .ZN(_04085_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09206_ (.A1(_04083_),
    .A2(_04084_),
    .B1(_04085_),
    .B2(_02589_),
    .ZN(_04086_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09207_ (.A1(_02557_),
    .A2(_04086_),
    .Z(_04087_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09208_ (.A1(_02703_),
    .A2(_04087_),
    .B(_00703_),
    .C(_02676_),
    .ZN(_04088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09209_ (.A1(_04078_),
    .A2(_04088_),
    .ZN(_00729_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09210_ (.A1(_04034_),
    .A2(_02628_),
    .A3(_00710_),
    .Z(_04089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09211_ (.I(_04089_),
    .Z(_00730_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09212_ (.A1(_02597_),
    .A2(_04038_),
    .ZN(_04090_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09213_ (.A1(_03112_),
    .A2(_04027_),
    .B(_04090_),
    .ZN(_00731_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09214_ (.I(_02730_),
    .Z(_04091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09215_ (.A1(_04091_),
    .A2(_02982_),
    .ZN(_04092_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09216_ (.I(_04092_),
    .Z(_04093_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09217_ (.I(_04092_),
    .Z(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09218_ (.A1(\u_cpu.rf_ram.memory[92][0] ),
    .A2(_04094_),
    .ZN(_04095_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09219_ (.A1(_04056_),
    .A2(_04093_),
    .B(_04095_),
    .ZN(_00732_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09220_ (.A1(\u_cpu.rf_ram.memory[92][1] ),
    .A2(_04094_),
    .ZN(_04096_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09221_ (.A1(_04061_),
    .A2(_04093_),
    .B(_04096_),
    .ZN(_00733_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09222_ (.I(_04092_),
    .Z(_04097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09223_ (.A1(\u_cpu.rf_ram.memory[92][2] ),
    .A2(_04097_),
    .ZN(_04098_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09224_ (.A1(_04063_),
    .A2(_04093_),
    .B(_04098_),
    .ZN(_00734_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09225_ (.A1(\u_cpu.rf_ram.memory[92][3] ),
    .A2(_04097_),
    .ZN(_04099_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09226_ (.A1(_04066_),
    .A2(_04093_),
    .B(_04099_),
    .ZN(_00735_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09227_ (.A1(\u_cpu.rf_ram.memory[92][4] ),
    .A2(_04097_),
    .ZN(_04100_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09228_ (.A1(_04068_),
    .A2(_04093_),
    .B(_04100_),
    .ZN(_00736_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09229_ (.A1(\u_cpu.rf_ram.memory[92][5] ),
    .A2(_04097_),
    .ZN(_04101_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09230_ (.A1(_04070_),
    .A2(_04094_),
    .B(_04101_),
    .ZN(_00737_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09231_ (.A1(\u_cpu.rf_ram.memory[92][6] ),
    .A2(_04097_),
    .ZN(_04102_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09232_ (.A1(_04072_),
    .A2(_04094_),
    .B(_04102_),
    .ZN(_00738_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09233_ (.A1(\u_cpu.rf_ram.memory[92][7] ),
    .A2(_04092_),
    .ZN(_04103_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09234_ (.A1(_04074_),
    .A2(_04094_),
    .B(_04103_),
    .ZN(_00739_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09235_ (.A1(_02939_),
    .A2(_03310_),
    .ZN(_04104_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09236_ (.I(_04104_),
    .Z(_04105_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09237_ (.I(_04104_),
    .Z(_04106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09238_ (.A1(\u_cpu.rf_ram.memory[35][0] ),
    .A2(_04106_),
    .ZN(_04107_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09239_ (.A1(_04056_),
    .A2(_04105_),
    .B(_04107_),
    .ZN(_00740_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09240_ (.A1(\u_cpu.rf_ram.memory[35][1] ),
    .A2(_04106_),
    .ZN(_04108_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09241_ (.A1(_04061_),
    .A2(_04105_),
    .B(_04108_),
    .ZN(_00741_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09242_ (.I(_04104_),
    .Z(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09243_ (.A1(\u_cpu.rf_ram.memory[35][2] ),
    .A2(_04109_),
    .ZN(_04110_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09244_ (.A1(_04063_),
    .A2(_04105_),
    .B(_04110_),
    .ZN(_00742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09245_ (.A1(\u_cpu.rf_ram.memory[35][3] ),
    .A2(_04109_),
    .ZN(_04111_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09246_ (.A1(_04066_),
    .A2(_04105_),
    .B(_04111_),
    .ZN(_00743_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09247_ (.A1(\u_cpu.rf_ram.memory[35][4] ),
    .A2(_04109_),
    .ZN(_04112_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09248_ (.A1(_04068_),
    .A2(_04105_),
    .B(_04112_),
    .ZN(_00744_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09249_ (.A1(\u_cpu.rf_ram.memory[35][5] ),
    .A2(_04109_),
    .ZN(_04113_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09250_ (.A1(_04070_),
    .A2(_04106_),
    .B(_04113_),
    .ZN(_00745_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09251_ (.A1(\u_cpu.rf_ram.memory[35][6] ),
    .A2(_04109_),
    .ZN(_04114_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09252_ (.A1(_04072_),
    .A2(_04106_),
    .B(_04114_),
    .ZN(_00746_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09253_ (.A1(\u_cpu.rf_ram.memory[35][7] ),
    .A2(_04104_),
    .ZN(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09254_ (.A1(_04074_),
    .A2(_04106_),
    .B(_04115_),
    .ZN(_00747_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09255_ (.A1(_02722_),
    .A2(_02965_),
    .ZN(_04116_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09256_ (.I(_04116_),
    .Z(_04117_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09257_ (.I(_04116_),
    .Z(_04118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09258_ (.A1(\u_cpu.rf_ram.memory[34][0] ),
    .A2(_04118_),
    .ZN(_04119_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09259_ (.A1(_04056_),
    .A2(_04117_),
    .B(_04119_),
    .ZN(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09260_ (.A1(\u_cpu.rf_ram.memory[34][1] ),
    .A2(_04118_),
    .ZN(_04120_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09261_ (.A1(_04061_),
    .A2(_04117_),
    .B(_04120_),
    .ZN(_00749_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09262_ (.I(_04116_),
    .Z(_04121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09263_ (.A1(\u_cpu.rf_ram.memory[34][2] ),
    .A2(_04121_),
    .ZN(_04122_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09264_ (.A1(_04063_),
    .A2(_04117_),
    .B(_04122_),
    .ZN(_00750_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09265_ (.A1(\u_cpu.rf_ram.memory[34][3] ),
    .A2(_04121_),
    .ZN(_04123_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09266_ (.A1(_04066_),
    .A2(_04117_),
    .B(_04123_),
    .ZN(_00751_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09267_ (.A1(\u_cpu.rf_ram.memory[34][4] ),
    .A2(_04121_),
    .ZN(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09268_ (.A1(_04068_),
    .A2(_04117_),
    .B(_04124_),
    .ZN(_00752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09269_ (.A1(\u_cpu.rf_ram.memory[34][5] ),
    .A2(_04121_),
    .ZN(_04125_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09270_ (.A1(_04070_),
    .A2(_04118_),
    .B(_04125_),
    .ZN(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09271_ (.A1(\u_cpu.rf_ram.memory[34][6] ),
    .A2(_04121_),
    .ZN(_04126_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09272_ (.A1(_04072_),
    .A2(_04118_),
    .B(_04126_),
    .ZN(_00754_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09273_ (.A1(\u_cpu.rf_ram.memory[34][7] ),
    .A2(_04116_),
    .ZN(_04127_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09274_ (.A1(_04074_),
    .A2(_04118_),
    .B(_04127_),
    .ZN(_00755_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09275_ (.A1(_02785_),
    .A2(_03970_),
    .ZN(_04128_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09276_ (.I(_04128_),
    .Z(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09277_ (.I(_04128_),
    .Z(_04130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09278_ (.A1(\u_cpu.rf_ram.memory[117][0] ),
    .A2(_04130_),
    .ZN(_04131_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09279_ (.A1(_04056_),
    .A2(_04129_),
    .B(_04131_),
    .ZN(_00756_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09280_ (.A1(\u_cpu.rf_ram.memory[117][1] ),
    .A2(_04130_),
    .ZN(_04132_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09281_ (.A1(_04061_),
    .A2(_04129_),
    .B(_04132_),
    .ZN(_00757_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09282_ (.I(_04128_),
    .Z(_04133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09283_ (.A1(\u_cpu.rf_ram.memory[117][2] ),
    .A2(_04133_),
    .ZN(_04134_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09284_ (.A1(_04063_),
    .A2(_04129_),
    .B(_04134_),
    .ZN(_00758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09285_ (.A1(\u_cpu.rf_ram.memory[117][3] ),
    .A2(_04133_),
    .ZN(_04135_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09286_ (.A1(_04066_),
    .A2(_04129_),
    .B(_04135_),
    .ZN(_00759_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09287_ (.A1(\u_cpu.rf_ram.memory[117][4] ),
    .A2(_04133_),
    .ZN(_04136_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09288_ (.A1(_04068_),
    .A2(_04129_),
    .B(_04136_),
    .ZN(_00760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09289_ (.A1(\u_cpu.rf_ram.memory[117][5] ),
    .A2(_04133_),
    .ZN(_04137_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09290_ (.A1(_04070_),
    .A2(_04130_),
    .B(_04137_),
    .ZN(_00761_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09291_ (.A1(\u_cpu.rf_ram.memory[117][6] ),
    .A2(_04133_),
    .ZN(_04138_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09292_ (.A1(_04072_),
    .A2(_04130_),
    .B(_04138_),
    .ZN(_00762_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09293_ (.A1(\u_cpu.rf_ram.memory[117][7] ),
    .A2(_04128_),
    .ZN(_04139_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09294_ (.A1(_04074_),
    .A2(_04130_),
    .B(_04139_),
    .ZN(_00763_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09295_ (.I(_03893_),
    .Z(_04140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09296_ (.A1(_03165_),
    .A2(_03970_),
    .ZN(_04141_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09297_ (.I(_04141_),
    .Z(_04142_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09298_ (.I(_04141_),
    .Z(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09299_ (.A1(\u_cpu.rf_ram.memory[120][0] ),
    .A2(_04143_),
    .ZN(_04144_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09300_ (.A1(_04140_),
    .A2(_04142_),
    .B(_04144_),
    .ZN(_00764_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09301_ (.I(_03899_),
    .Z(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09302_ (.A1(\u_cpu.rf_ram.memory[120][1] ),
    .A2(_04143_),
    .ZN(_04146_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09303_ (.A1(_04145_),
    .A2(_04142_),
    .B(_04146_),
    .ZN(_00765_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09304_ (.I(_03902_),
    .Z(_04147_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09305_ (.I(_04141_),
    .Z(_04148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09306_ (.A1(\u_cpu.rf_ram.memory[120][2] ),
    .A2(_04148_),
    .ZN(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09307_ (.A1(_04147_),
    .A2(_04142_),
    .B(_04149_),
    .ZN(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09308_ (.I(_03906_),
    .Z(_04150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09309_ (.A1(\u_cpu.rf_ram.memory[120][3] ),
    .A2(_04148_),
    .ZN(_04151_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09310_ (.A1(_04150_),
    .A2(_04142_),
    .B(_04151_),
    .ZN(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09311_ (.I(_03909_),
    .Z(_04152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09312_ (.A1(\u_cpu.rf_ram.memory[120][4] ),
    .A2(_04148_),
    .ZN(_04153_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09313_ (.A1(_04152_),
    .A2(_04142_),
    .B(_04153_),
    .ZN(_00768_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09314_ (.I(_03912_),
    .Z(_04154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09315_ (.A1(\u_cpu.rf_ram.memory[120][5] ),
    .A2(_04148_),
    .ZN(_04155_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09316_ (.A1(_04154_),
    .A2(_04143_),
    .B(_04155_),
    .ZN(_00769_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09317_ (.I(_03915_),
    .Z(_04156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09318_ (.A1(\u_cpu.rf_ram.memory[120][6] ),
    .A2(_04148_),
    .ZN(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09319_ (.A1(_04156_),
    .A2(_04143_),
    .B(_04157_),
    .ZN(_00770_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09320_ (.I(_03918_),
    .Z(_04158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09321_ (.A1(\u_cpu.rf_ram.memory[120][7] ),
    .A2(_04141_),
    .ZN(_04159_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09322_ (.A1(_04158_),
    .A2(_04143_),
    .B(_04159_),
    .ZN(_00771_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09323_ (.A1(_03180_),
    .A2(_03286_),
    .ZN(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09324_ (.I(_04160_),
    .Z(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09325_ (.I(_04160_),
    .Z(_04162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09326_ (.A1(\u_cpu.rf_ram.memory[118][0] ),
    .A2(_04162_),
    .ZN(_04163_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09327_ (.A1(_04140_),
    .A2(_04161_),
    .B(_04163_),
    .ZN(_00772_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09328_ (.A1(\u_cpu.rf_ram.memory[118][1] ),
    .A2(_04162_),
    .ZN(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09329_ (.A1(_04145_),
    .A2(_04161_),
    .B(_04164_),
    .ZN(_00773_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09330_ (.I(_04160_),
    .Z(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09331_ (.A1(\u_cpu.rf_ram.memory[118][2] ),
    .A2(_04165_),
    .ZN(_04166_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09332_ (.A1(_04147_),
    .A2(_04161_),
    .B(_04166_),
    .ZN(_00774_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09333_ (.A1(\u_cpu.rf_ram.memory[118][3] ),
    .A2(_04165_),
    .ZN(_04167_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09334_ (.A1(_04150_),
    .A2(_04161_),
    .B(_04167_),
    .ZN(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09335_ (.A1(\u_cpu.rf_ram.memory[118][4] ),
    .A2(_04165_),
    .ZN(_04168_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09336_ (.A1(_04152_),
    .A2(_04161_),
    .B(_04168_),
    .ZN(_00776_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09337_ (.A1(\u_cpu.rf_ram.memory[118][5] ),
    .A2(_04165_),
    .ZN(_04169_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09338_ (.A1(_04154_),
    .A2(_04162_),
    .B(_04169_),
    .ZN(_00777_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09339_ (.A1(\u_cpu.rf_ram.memory[118][6] ),
    .A2(_04165_),
    .ZN(_04170_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09340_ (.A1(_04156_),
    .A2(_04162_),
    .B(_04170_),
    .ZN(_00778_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09341_ (.A1(\u_cpu.rf_ram.memory[118][7] ),
    .A2(_04160_),
    .ZN(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09342_ (.A1(_04158_),
    .A2(_04162_),
    .B(_04171_),
    .ZN(_00779_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09343_ (.A1(_03019_),
    .A2(_03970_),
    .ZN(_04172_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09344_ (.I(_04172_),
    .Z(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09345_ (.I(_04172_),
    .Z(_04174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09346_ (.A1(\u_cpu.rf_ram.memory[121][0] ),
    .A2(_04174_),
    .ZN(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09347_ (.A1(_04140_),
    .A2(_04173_),
    .B(_04175_),
    .ZN(_00780_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09348_ (.A1(\u_cpu.rf_ram.memory[121][1] ),
    .A2(_04174_),
    .ZN(_04176_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09349_ (.A1(_04145_),
    .A2(_04173_),
    .B(_04176_),
    .ZN(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09350_ (.I(_04172_),
    .Z(_04177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09351_ (.A1(\u_cpu.rf_ram.memory[121][2] ),
    .A2(_04177_),
    .ZN(_04178_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09352_ (.A1(_04147_),
    .A2(_04173_),
    .B(_04178_),
    .ZN(_00782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09353_ (.A1(\u_cpu.rf_ram.memory[121][3] ),
    .A2(_04177_),
    .ZN(_04179_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09354_ (.A1(_04150_),
    .A2(_04173_),
    .B(_04179_),
    .ZN(_00783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09355_ (.A1(\u_cpu.rf_ram.memory[121][4] ),
    .A2(_04177_),
    .ZN(_04180_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09356_ (.A1(_04152_),
    .A2(_04173_),
    .B(_04180_),
    .ZN(_00784_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09357_ (.A1(\u_cpu.rf_ram.memory[121][5] ),
    .A2(_04177_),
    .ZN(_04181_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09358_ (.A1(_04154_),
    .A2(_04174_),
    .B(_04181_),
    .ZN(_00785_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09359_ (.A1(\u_cpu.rf_ram.memory[121][6] ),
    .A2(_04177_),
    .ZN(_04182_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09360_ (.A1(_04156_),
    .A2(_04174_),
    .B(_04182_),
    .ZN(_00786_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09361_ (.A1(\u_cpu.rf_ram.memory[121][7] ),
    .A2(_04172_),
    .ZN(_04183_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09362_ (.A1(_04158_),
    .A2(_04174_),
    .B(_04183_),
    .ZN(_00787_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09363_ (.I(_02845_),
    .Z(_04184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09364_ (.A1(_03870_),
    .A2(_03166_),
    .ZN(_04185_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09365_ (.I(_04185_),
    .Z(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09366_ (.I0(_04184_),
    .I1(\u_cpu.rf_ram.memory[8][0] ),
    .S(_04186_),
    .Z(_04187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09367_ (.I(_04187_),
    .Z(_00788_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09368_ (.I(_02854_),
    .Z(_04188_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09369_ (.I0(_04188_),
    .I1(\u_cpu.rf_ram.memory[8][1] ),
    .S(_04186_),
    .Z(_04189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09370_ (.I(_04189_),
    .Z(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09371_ (.I(_02857_),
    .Z(_04190_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09372_ (.I0(_04190_),
    .I1(\u_cpu.rf_ram.memory[8][2] ),
    .S(_04186_),
    .Z(_04191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09373_ (.I(_04191_),
    .Z(_00790_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09374_ (.I(_02860_),
    .Z(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09375_ (.I0(_04192_),
    .I1(\u_cpu.rf_ram.memory[8][3] ),
    .S(_04186_),
    .Z(_04193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09376_ (.I(_04193_),
    .Z(_00791_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09377_ (.I(_02863_),
    .Z(_04194_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09378_ (.I0(_04194_),
    .I1(\u_cpu.rf_ram.memory[8][4] ),
    .S(_04186_),
    .Z(_04195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09379_ (.I(_04195_),
    .Z(_00792_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09380_ (.I(_02866_),
    .Z(_04196_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09381_ (.I0(_04196_),
    .I1(\u_cpu.rf_ram.memory[8][5] ),
    .S(_04185_),
    .Z(_04197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09382_ (.I(_04197_),
    .Z(_00793_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09383_ (.I(_02869_),
    .Z(_04198_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09384_ (.I0(_04198_),
    .I1(\u_cpu.rf_ram.memory[8][6] ),
    .S(_04185_),
    .Z(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09385_ (.I(_04199_),
    .Z(_00794_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09386_ (.I(_02872_),
    .Z(_04200_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09387_ (.I0(_04200_),
    .I1(\u_cpu.rf_ram.memory[8][7] ),
    .S(_04185_),
    .Z(_04201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09388_ (.I(_04201_),
    .Z(_00795_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09389_ (.A1(_03870_),
    .A2(_03034_),
    .ZN(_04202_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09390_ (.I(_04202_),
    .Z(_04203_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09391_ (.I0(_04184_),
    .I1(\u_cpu.rf_ram.memory[11][0] ),
    .S(_04203_),
    .Z(_04204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09392_ (.I(_04204_),
    .Z(_00796_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09393_ (.I0(_04188_),
    .I1(\u_cpu.rf_ram.memory[11][1] ),
    .S(_04203_),
    .Z(_04205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09394_ (.I(_04205_),
    .Z(_00797_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09395_ (.I0(_04190_),
    .I1(\u_cpu.rf_ram.memory[11][2] ),
    .S(_04203_),
    .Z(_04206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09396_ (.I(_04206_),
    .Z(_00798_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09397_ (.I0(_04192_),
    .I1(\u_cpu.rf_ram.memory[11][3] ),
    .S(_04203_),
    .Z(_04207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09398_ (.I(_04207_),
    .Z(_00799_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09399_ (.I0(_04194_),
    .I1(\u_cpu.rf_ram.memory[11][4] ),
    .S(_04203_),
    .Z(_04208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09400_ (.I(_04208_),
    .Z(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09401_ (.I0(_04196_),
    .I1(\u_cpu.rf_ram.memory[11][5] ),
    .S(_04202_),
    .Z(_04209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09402_ (.I(_04209_),
    .Z(_00801_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09403_ (.I0(_04198_),
    .I1(\u_cpu.rf_ram.memory[11][6] ),
    .S(_04202_),
    .Z(_04210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09404_ (.I(_04210_),
    .Z(_00802_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09405_ (.I0(_04200_),
    .I1(\u_cpu.rf_ram.memory[11][7] ),
    .S(_04202_),
    .Z(_04211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09406_ (.I(_04211_),
    .Z(_00803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09407_ (.A1(_02890_),
    .A2(_03970_),
    .ZN(_04212_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09408_ (.I(_04212_),
    .Z(_04213_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09409_ (.I(_04212_),
    .Z(_04214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09410_ (.A1(\u_cpu.rf_ram.memory[112][0] ),
    .A2(_04214_),
    .ZN(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09411_ (.A1(_04140_),
    .A2(_04213_),
    .B(_04215_),
    .ZN(_00804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09412_ (.A1(\u_cpu.rf_ram.memory[112][1] ),
    .A2(_04214_),
    .ZN(_04216_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09413_ (.A1(_04145_),
    .A2(_04213_),
    .B(_04216_),
    .ZN(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09414_ (.I(_04212_),
    .Z(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09415_ (.A1(\u_cpu.rf_ram.memory[112][2] ),
    .A2(_04217_),
    .ZN(_04218_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09416_ (.A1(_04147_),
    .A2(_04213_),
    .B(_04218_),
    .ZN(_00806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09417_ (.A1(\u_cpu.rf_ram.memory[112][3] ),
    .A2(_04217_),
    .ZN(_04219_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09418_ (.A1(_04150_),
    .A2(_04213_),
    .B(_04219_),
    .ZN(_00807_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09419_ (.A1(\u_cpu.rf_ram.memory[112][4] ),
    .A2(_04217_),
    .ZN(_04220_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09420_ (.A1(_04152_),
    .A2(_04213_),
    .B(_04220_),
    .ZN(_00808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09421_ (.A1(\u_cpu.rf_ram.memory[112][5] ),
    .A2(_04217_),
    .ZN(_04221_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09422_ (.A1(_04154_),
    .A2(_04214_),
    .B(_04221_),
    .ZN(_00809_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09423_ (.A1(\u_cpu.rf_ram.memory[112][6] ),
    .A2(_04217_),
    .ZN(_04222_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09424_ (.A1(_04156_),
    .A2(_04214_),
    .B(_04222_),
    .ZN(_00810_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09425_ (.A1(\u_cpu.rf_ram.memory[112][7] ),
    .A2(_04212_),
    .ZN(_04223_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09426_ (.A1(_04158_),
    .A2(_04214_),
    .B(_04223_),
    .ZN(_00811_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09427_ (.I(_03180_),
    .Z(_04224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09428_ (.A1(_02937_),
    .A2(_04224_),
    .ZN(_04225_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09429_ (.I(_04225_),
    .Z(_04226_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09430_ (.I(_04225_),
    .Z(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09431_ (.A1(\u_cpu.rf_ram.memory[122][0] ),
    .A2(_04227_),
    .ZN(_04228_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09432_ (.A1(_04140_),
    .A2(_04226_),
    .B(_04228_),
    .ZN(_00812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09433_ (.A1(\u_cpu.rf_ram.memory[122][1] ),
    .A2(_04227_),
    .ZN(_04229_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09434_ (.A1(_04145_),
    .A2(_04226_),
    .B(_04229_),
    .ZN(_00813_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09435_ (.I(_04225_),
    .Z(_04230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09436_ (.A1(\u_cpu.rf_ram.memory[122][2] ),
    .A2(_04230_),
    .ZN(_04231_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09437_ (.A1(_04147_),
    .A2(_04226_),
    .B(_04231_),
    .ZN(_00814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09438_ (.A1(\u_cpu.rf_ram.memory[122][3] ),
    .A2(_04230_),
    .ZN(_04232_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09439_ (.A1(_04150_),
    .A2(_04226_),
    .B(_04232_),
    .ZN(_00815_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09440_ (.A1(\u_cpu.rf_ram.memory[122][4] ),
    .A2(_04230_),
    .ZN(_04233_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09441_ (.A1(_04152_),
    .A2(_04226_),
    .B(_04233_),
    .ZN(_00816_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09442_ (.A1(\u_cpu.rf_ram.memory[122][5] ),
    .A2(_04230_),
    .ZN(_04234_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09443_ (.A1(_04154_),
    .A2(_04227_),
    .B(_04234_),
    .ZN(_00817_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09444_ (.A1(\u_cpu.rf_ram.memory[122][6] ),
    .A2(_04230_),
    .ZN(_04235_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09445_ (.A1(_04156_),
    .A2(_04227_),
    .B(_04235_),
    .ZN(_00818_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09446_ (.A1(\u_cpu.rf_ram.memory[122][7] ),
    .A2(_04225_),
    .ZN(_04236_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09447_ (.A1(_04158_),
    .A2(_04227_),
    .B(_04236_),
    .ZN(_00819_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09448_ (.I(_03893_),
    .Z(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09449_ (.A1(_03002_),
    .A2(_04224_),
    .ZN(_04238_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09450_ (.I(_04238_),
    .Z(_04239_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09451_ (.I(_04238_),
    .Z(_04240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09452_ (.A1(\u_cpu.rf_ram.memory[115][0] ),
    .A2(_04240_),
    .ZN(_04241_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09453_ (.A1(_04237_),
    .A2(_04239_),
    .B(_04241_),
    .ZN(_00820_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09454_ (.I(_03899_),
    .Z(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09455_ (.A1(\u_cpu.rf_ram.memory[115][1] ),
    .A2(_04240_),
    .ZN(_04243_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09456_ (.A1(_04242_),
    .A2(_04239_),
    .B(_04243_),
    .ZN(_00821_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09457_ (.I(_03902_),
    .Z(_04244_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09458_ (.I(_04238_),
    .Z(_04245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09459_ (.A1(\u_cpu.rf_ram.memory[115][2] ),
    .A2(_04245_),
    .ZN(_04246_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09460_ (.A1(_04244_),
    .A2(_04239_),
    .B(_04246_),
    .ZN(_00822_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09461_ (.I(_03906_),
    .Z(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09462_ (.A1(\u_cpu.rf_ram.memory[115][3] ),
    .A2(_04245_),
    .ZN(_04248_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09463_ (.A1(_04247_),
    .A2(_04239_),
    .B(_04248_),
    .ZN(_00823_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09464_ (.I(_03909_),
    .Z(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09465_ (.A1(\u_cpu.rf_ram.memory[115][4] ),
    .A2(_04245_),
    .ZN(_04250_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09466_ (.A1(_04249_),
    .A2(_04239_),
    .B(_04250_),
    .ZN(_00824_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09467_ (.I(_03912_),
    .Z(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09468_ (.A1(\u_cpu.rf_ram.memory[115][5] ),
    .A2(_04245_),
    .ZN(_04252_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09469_ (.A1(_04251_),
    .A2(_04240_),
    .B(_04252_),
    .ZN(_00825_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09470_ (.I(_03915_),
    .Z(_04253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09471_ (.A1(\u_cpu.rf_ram.memory[115][6] ),
    .A2(_04245_),
    .ZN(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09472_ (.A1(_04253_),
    .A2(_04240_),
    .B(_04254_),
    .ZN(_00826_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09473_ (.I(_03918_),
    .Z(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09474_ (.A1(\u_cpu.rf_ram.memory[115][7] ),
    .A2(_04238_),
    .ZN(_04256_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09475_ (.A1(_04255_),
    .A2(_04240_),
    .B(_04256_),
    .ZN(_00827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09476_ (.A1(_02830_),
    .A2(_04224_),
    .ZN(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09477_ (.I(_04257_),
    .Z(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09478_ (.I(_04257_),
    .Z(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09479_ (.A1(\u_cpu.rf_ram.memory[116][0] ),
    .A2(_04259_),
    .ZN(_04260_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09480_ (.A1(_04237_),
    .A2(_04258_),
    .B(_04260_),
    .ZN(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09481_ (.A1(\u_cpu.rf_ram.memory[116][1] ),
    .A2(_04259_),
    .ZN(_04261_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09482_ (.A1(_04242_),
    .A2(_04258_),
    .B(_04261_),
    .ZN(_00829_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09483_ (.I(_04257_),
    .Z(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09484_ (.A1(\u_cpu.rf_ram.memory[116][2] ),
    .A2(_04262_),
    .ZN(_04263_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09485_ (.A1(_04244_),
    .A2(_04258_),
    .B(_04263_),
    .ZN(_00830_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09486_ (.A1(\u_cpu.rf_ram.memory[116][3] ),
    .A2(_04262_),
    .ZN(_04264_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09487_ (.A1(_04247_),
    .A2(_04258_),
    .B(_04264_),
    .ZN(_00831_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09488_ (.A1(\u_cpu.rf_ram.memory[116][4] ),
    .A2(_04262_),
    .ZN(_04265_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09489_ (.A1(_04249_),
    .A2(_04258_),
    .B(_04265_),
    .ZN(_00832_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09490_ (.A1(\u_cpu.rf_ram.memory[116][5] ),
    .A2(_04262_),
    .ZN(_04266_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09491_ (.A1(_04251_),
    .A2(_04259_),
    .B(_04266_),
    .ZN(_00833_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09492_ (.A1(\u_cpu.rf_ram.memory[116][6] ),
    .A2(_04262_),
    .ZN(_04267_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09493_ (.A1(_04253_),
    .A2(_04259_),
    .B(_04267_),
    .ZN(_00834_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09494_ (.A1(\u_cpu.rf_ram.memory[116][7] ),
    .A2(_04257_),
    .ZN(_04268_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09495_ (.A1(_04255_),
    .A2(_04259_),
    .B(_04268_),
    .ZN(_00835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09496_ (.A1(_02803_),
    .A2(_02965_),
    .ZN(_04269_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09497_ (.I(_04269_),
    .Z(_04270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09498_ (.I(_04269_),
    .Z(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09499_ (.A1(\u_cpu.rf_ram.memory[33][0] ),
    .A2(_04271_),
    .ZN(_04272_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09500_ (.A1(_04237_),
    .A2(_04270_),
    .B(_04272_),
    .ZN(_00836_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09501_ (.A1(\u_cpu.rf_ram.memory[33][1] ),
    .A2(_04271_),
    .ZN(_04273_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09502_ (.A1(_04242_),
    .A2(_04270_),
    .B(_04273_),
    .ZN(_00837_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09503_ (.I(_04269_),
    .Z(_04274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09504_ (.A1(\u_cpu.rf_ram.memory[33][2] ),
    .A2(_04274_),
    .ZN(_04275_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09505_ (.A1(_04244_),
    .A2(_04270_),
    .B(_04275_),
    .ZN(_00838_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09506_ (.A1(\u_cpu.rf_ram.memory[33][3] ),
    .A2(_04274_),
    .ZN(_04276_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09507_ (.A1(_04247_),
    .A2(_04270_),
    .B(_04276_),
    .ZN(_00839_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09508_ (.A1(\u_cpu.rf_ram.memory[33][4] ),
    .A2(_04274_),
    .ZN(_04277_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09509_ (.A1(_04249_),
    .A2(_04270_),
    .B(_04277_),
    .ZN(_00840_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09510_ (.A1(\u_cpu.rf_ram.memory[33][5] ),
    .A2(_04274_),
    .ZN(_04278_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09511_ (.A1(_04251_),
    .A2(_04271_),
    .B(_04278_),
    .ZN(_00841_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09512_ (.A1(\u_cpu.rf_ram.memory[33][6] ),
    .A2(_04274_),
    .ZN(_04279_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09513_ (.A1(_04253_),
    .A2(_04271_),
    .B(_04279_),
    .ZN(_00842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09514_ (.A1(\u_cpu.rf_ram.memory[33][7] ),
    .A2(_04269_),
    .ZN(_04280_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09515_ (.A1(_04255_),
    .A2(_04271_),
    .B(_04280_),
    .ZN(_00843_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09516_ (.A1(\u_cpu.cpu.bufreg.lsb[1] ),
    .A2(_04034_),
    .B(_04031_),
    .C(_01369_),
    .ZN(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09517_ (.A1(_01370_),
    .A2(_04034_),
    .ZN(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09518_ (.A1(_02528_),
    .A2(_04281_),
    .A3(_04282_),
    .ZN(_04283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09519_ (.A1(_03122_),
    .A2(_04283_),
    .ZN(_04284_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09520_ (.I(_04284_),
    .Z(_04285_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09521_ (.I(_03124_),
    .Z(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09522_ (.A1(_03125_),
    .A2(_04286_),
    .ZN(_04287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09523_ (.A1(_04285_),
    .A2(_04287_),
    .ZN(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09524_ (.I(_03124_),
    .Z(_04289_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09525_ (.I(_03132_),
    .Z(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09526_ (.A1(net36),
    .A2(_04289_),
    .B(_04290_),
    .ZN(_04291_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09527_ (.A1(net8),
    .A2(_01450_),
    .Z(_04292_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09528_ (.I(_04292_),
    .Z(_04293_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09529_ (.A1(_04292_),
    .A2(_04284_),
    .ZN(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09530_ (.I(_04294_),
    .Z(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09531_ (.A1(\u_arbiter.i_wb_cpu_rdt[0] ),
    .A2(_04293_),
    .B1(_04295_),
    .B2(_03125_),
    .ZN(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09532_ (.A1(_04288_),
    .A2(_04291_),
    .B(_04296_),
    .ZN(_00844_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09533_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[2] ),
    .A2(_04286_),
    .ZN(_04297_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09534_ (.A1(_03125_),
    .A2(net36),
    .B(_04286_),
    .ZN(_04298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09535_ (.A1(_04285_),
    .A2(_04298_),
    .ZN(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09536_ (.I(_03132_),
    .Z(_04300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09537_ (.A1(net36),
    .A2(_04288_),
    .ZN(_04301_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09538_ (.A1(_04297_),
    .A2(_04299_),
    .B(_04300_),
    .C(_04301_),
    .ZN(_04302_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09539_ (.A1(\u_arbiter.i_wb_cpu_rdt[1] ),
    .A2(_04290_),
    .B(_04302_),
    .ZN(_04303_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09540_ (.I(_04303_),
    .ZN(_00845_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09541_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[3] ),
    .A2(_04286_),
    .ZN(_04304_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09542_ (.A1(_03125_),
    .A2(net36),
    .A3(\u_arbiter.i_wb_cpu_dbus_dat[2] ),
    .B(_04286_),
    .ZN(_04305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09543_ (.A1(_04285_),
    .A2(_04305_),
    .ZN(_04306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09544_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[2] ),
    .A2(_04299_),
    .ZN(_04307_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09545_ (.A1(_04304_),
    .A2(_04306_),
    .B(_04300_),
    .C(_04307_),
    .ZN(_04308_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09546_ (.A1(\u_arbiter.i_wb_cpu_rdt[2] ),
    .A2(_04290_),
    .B(_04308_),
    .ZN(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09547_ (.I(_04309_),
    .ZN(_00846_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _09548_ (.I(\u_arbiter.i_wb_cpu_rdt[3] ),
    .ZN(_04310_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09549_ (.I(_04292_),
    .Z(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09550_ (.I(_04311_),
    .Z(_04312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09551_ (.A1(_04289_),
    .A2(_03126_),
    .ZN(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09552_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[4] ),
    .A2(_04289_),
    .B(_04285_),
    .C(_04313_),
    .ZN(_04314_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09553_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[3] ),
    .A2(_04306_),
    .B(_04311_),
    .ZN(_04315_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09554_ (.A1(_04310_),
    .A2(_04312_),
    .B1(_04314_),
    .B2(_04315_),
    .ZN(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09555_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[4] ),
    .A2(_03126_),
    .Z(_04316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09556_ (.A1(_04289_),
    .A2(_04316_),
    .ZN(_04317_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09557_ (.A1(_03132_),
    .A2(_04284_),
    .Z(_04318_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09558_ (.I(_04318_),
    .Z(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09559_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .A2(_04289_),
    .B(_04317_),
    .C(_04319_),
    .ZN(_04320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09560_ (.I(_04294_),
    .Z(_04321_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09561_ (.I(_04321_),
    .Z(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09562_ (.A1(\u_arbiter.i_wb_cpu_rdt[4] ),
    .A2(_04312_),
    .B1(_04322_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[4] ),
    .ZN(_04323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09563_ (.A1(_04320_),
    .A2(_04323_),
    .ZN(_00848_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09564_ (.A1(\u_arbiter.i_wb_cpu_rdt[5] ),
    .A2(_04312_),
    .ZN(_04324_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09565_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .A2(_04295_),
    .B1(_04319_),
    .B2(_03130_),
    .ZN(_04325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09566_ (.A1(_04324_),
    .A2(_04325_),
    .ZN(_00849_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09567_ (.I(_04292_),
    .Z(_04326_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09568_ (.I(_04318_),
    .Z(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _09569_ (.A1(\u_arbiter.i_wb_cpu_rdt[6] ),
    .A2(_04326_),
    .B1(_04321_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[6] ),
    .C1(_04327_),
    .C2(\u_arbiter.i_wb_cpu_dbus_dat[7] ),
    .ZN(_04328_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09570_ (.I(_04328_),
    .ZN(_00850_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09571_ (.I(_04327_),
    .Z(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09572_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[8] ),
    .A2(_04329_),
    .ZN(_04330_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09573_ (.I(_04294_),
    .Z(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09574_ (.A1(\u_arbiter.i_wb_cpu_rdt[7] ),
    .A2(_04312_),
    .B1(_04331_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[7] ),
    .ZN(_04332_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09575_ (.A1(_04330_),
    .A2(_04332_),
    .ZN(_00851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09576_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[9] ),
    .A2(_04329_),
    .ZN(_04333_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09577_ (.I(_04311_),
    .Z(_04334_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09578_ (.A1(\u_arbiter.i_wb_cpu_rdt[8] ),
    .A2(_04334_),
    .B1(_04331_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[8] ),
    .ZN(_04335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09579_ (.A1(_04333_),
    .A2(_04335_),
    .ZN(_00852_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09580_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[10] ),
    .A2(_04329_),
    .ZN(_04336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09581_ (.A1(\u_arbiter.i_wb_cpu_rdt[9] ),
    .A2(_04334_),
    .B1(_04331_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[9] ),
    .ZN(_04337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09582_ (.A1(_04336_),
    .A2(_04337_),
    .ZN(_00853_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09583_ (.I(_04318_),
    .Z(_04338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09584_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[11] ),
    .A2(_04338_),
    .ZN(_04339_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09585_ (.A1(\u_arbiter.i_wb_cpu_rdt[10] ),
    .A2(_04334_),
    .B1(_04331_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[10] ),
    .ZN(_04340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09586_ (.A1(_04339_),
    .A2(_04340_),
    .ZN(_00854_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09587_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[12] ),
    .A2(_04338_),
    .ZN(_04341_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09588_ (.A1(\u_arbiter.i_wb_cpu_rdt[11] ),
    .A2(_04334_),
    .B1(_04331_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[11] ),
    .ZN(_04342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09589_ (.A1(_04341_),
    .A2(_04342_),
    .ZN(_00855_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09590_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[13] ),
    .A2(_04338_),
    .ZN(_04343_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09591_ (.I(_04294_),
    .Z(_04344_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09592_ (.A1(\u_arbiter.i_wb_cpu_rdt[12] ),
    .A2(_04334_),
    .B1(_04344_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[12] ),
    .ZN(_04345_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09593_ (.A1(_04343_),
    .A2(_04345_),
    .ZN(_00856_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09594_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[14] ),
    .A2(_04338_),
    .ZN(_04346_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09595_ (.I(_04311_),
    .Z(_04347_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09596_ (.A1(\u_arbiter.i_wb_cpu_rdt[13] ),
    .A2(_04347_),
    .B1(_04344_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[13] ),
    .ZN(_04348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09597_ (.A1(_04346_),
    .A2(_04348_),
    .ZN(_00857_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _09598_ (.A1(\u_arbiter.i_wb_cpu_rdt[14] ),
    .A2(_04326_),
    .B1(_04321_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[14] ),
    .C1(_04327_),
    .C2(\u_arbiter.i_wb_cpu_dbus_dat[15] ),
    .ZN(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09599_ (.I(_04349_),
    .ZN(_00858_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09600_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[16] ),
    .A2(_04338_),
    .ZN(_04350_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09601_ (.A1(\u_arbiter.i_wb_cpu_rdt[15] ),
    .A2(_04347_),
    .B1(_04344_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[15] ),
    .ZN(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09602_ (.A1(_04350_),
    .A2(_04351_),
    .ZN(_00859_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09603_ (.I(_04318_),
    .Z(_04352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09604_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[17] ),
    .A2(_04352_),
    .ZN(_04353_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09605_ (.A1(\u_arbiter.i_wb_cpu_rdt[16] ),
    .A2(_04347_),
    .B1(_04344_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[16] ),
    .ZN(_04354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09606_ (.A1(_04353_),
    .A2(_04354_),
    .ZN(_00860_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _09607_ (.A1(\u_arbiter.i_wb_cpu_rdt[17] ),
    .A2(_04326_),
    .B1(_04321_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[17] ),
    .C1(_04327_),
    .C2(\u_arbiter.i_wb_cpu_dbus_dat[18] ),
    .ZN(_04355_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09608_ (.I(_04355_),
    .ZN(_00861_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09609_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[19] ),
    .A2(_04352_),
    .ZN(_04356_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09610_ (.A1(\u_arbiter.i_wb_cpu_rdt[18] ),
    .A2(_04347_),
    .B1(_04344_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[18] ),
    .ZN(_04357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09611_ (.A1(_04356_),
    .A2(_04357_),
    .ZN(_00862_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09612_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[20] ),
    .A2(_04352_),
    .ZN(_04358_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09613_ (.I(_04294_),
    .Z(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09614_ (.A1(\u_arbiter.i_wb_cpu_rdt[19] ),
    .A2(_04347_),
    .B1(_04359_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[19] ),
    .ZN(_04360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09615_ (.A1(_04358_),
    .A2(_04360_),
    .ZN(_00863_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09616_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[21] ),
    .A2(_04352_),
    .ZN(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09617_ (.A1(\u_arbiter.i_wb_cpu_rdt[20] ),
    .A2(_04293_),
    .B1(_04359_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[20] ),
    .ZN(_04362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09618_ (.A1(_04361_),
    .A2(_04362_),
    .ZN(_00864_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _09619_ (.A1(\u_arbiter.i_wb_cpu_rdt[21] ),
    .A2(_04311_),
    .B1(_04321_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[21] ),
    .C1(_04327_),
    .C2(\u_arbiter.i_wb_cpu_dbus_dat[22] ),
    .ZN(_04363_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09620_ (.I(_04363_),
    .ZN(_00865_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09621_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[23] ),
    .A2(_04352_),
    .ZN(_04364_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09622_ (.A1(\u_arbiter.i_wb_cpu_rdt[22] ),
    .A2(_04293_),
    .B1(_04359_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[22] ),
    .ZN(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09623_ (.A1(_04364_),
    .A2(_04365_),
    .ZN(_00866_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09624_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[24] ),
    .A2(_04319_),
    .ZN(_04366_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09625_ (.A1(\u_arbiter.i_wb_cpu_rdt[23] ),
    .A2(_04293_),
    .B1(_04359_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[23] ),
    .ZN(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09626_ (.A1(_04366_),
    .A2(_04367_),
    .ZN(_00867_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09627_ (.A1(\u_arbiter.i_wb_cpu_rdt[24] ),
    .A2(_04312_),
    .ZN(_04368_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09628_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[24] ),
    .A2(_04295_),
    .B1(_04319_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[25] ),
    .ZN(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09629_ (.A1(_04368_),
    .A2(_04369_),
    .ZN(_00868_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09630_ (.I(\u_arbiter.i_wb_cpu_dbus_dat[26] ),
    .ZN(_04370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09631_ (.A1(_04300_),
    .A2(_04285_),
    .ZN(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09632_ (.A1(\u_arbiter.i_wb_cpu_rdt[25] ),
    .A2(_04326_),
    .B1(_04295_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[25] ),
    .ZN(_04372_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09633_ (.A1(_04370_),
    .A2(_04371_),
    .B(_04372_),
    .ZN(_00869_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09634_ (.A1(\u_arbiter.i_wb_cpu_rdt[26] ),
    .A2(_04290_),
    .B1(_04371_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[27] ),
    .ZN(_04373_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09635_ (.A1(_04370_),
    .A2(_04322_),
    .B(_04373_),
    .ZN(_00870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09636_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[28] ),
    .A2(_04319_),
    .ZN(_04374_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09637_ (.A1(\u_arbiter.i_wb_cpu_rdt[27] ),
    .A2(_04293_),
    .B1(_04359_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[27] ),
    .ZN(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09638_ (.A1(_04374_),
    .A2(_04375_),
    .ZN(_00871_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09639_ (.I(\u_arbiter.i_wb_cpu_dbus_dat[29] ),
    .ZN(_04376_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09640_ (.A1(\u_arbiter.i_wb_cpu_rdt[28] ),
    .A2(_04326_),
    .B1(_04295_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[28] ),
    .ZN(_04377_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09641_ (.A1(_04376_),
    .A2(_04371_),
    .B(_04377_),
    .ZN(_00872_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09642_ (.I(\u_arbiter.i_wb_cpu_dbus_dat[30] ),
    .ZN(_04378_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09643_ (.A1(\u_arbiter.i_wb_cpu_rdt[29] ),
    .A2(_04300_),
    .ZN(_04379_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09644_ (.A1(_04376_),
    .A2(_04322_),
    .B1(_04329_),
    .B2(_04378_),
    .C(_04379_),
    .ZN(_00873_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09645_ (.I(\u_arbiter.i_wb_cpu_dbus_dat[31] ),
    .ZN(_04380_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09646_ (.A1(\u_arbiter.i_wb_cpu_rdt[30] ),
    .A2(_04300_),
    .ZN(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09647_ (.A1(_04378_),
    .A2(_04322_),
    .B1(_04329_),
    .B2(_04380_),
    .C(_04381_),
    .ZN(_00874_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09648_ (.A1(\u_arbiter.i_wb_cpu_rdt[31] ),
    .A2(_04290_),
    .B1(_04371_),
    .B2(_02547_),
    .ZN(_04382_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09649_ (.A1(_04380_),
    .A2(_04322_),
    .B(_04382_),
    .ZN(_00875_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09650_ (.A1(_02803_),
    .A2(_04224_),
    .ZN(_04383_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09651_ (.I(_04383_),
    .Z(_04384_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09652_ (.I(_04383_),
    .Z(_04385_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09653_ (.A1(\u_cpu.rf_ram.memory[113][0] ),
    .A2(_04385_),
    .ZN(_04386_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09654_ (.A1(_04237_),
    .A2(_04384_),
    .B(_04386_),
    .ZN(_00876_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09655_ (.A1(\u_cpu.rf_ram.memory[113][1] ),
    .A2(_04385_),
    .ZN(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09656_ (.A1(_04242_),
    .A2(_04384_),
    .B(_04387_),
    .ZN(_00877_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09657_ (.I(_04383_),
    .Z(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09658_ (.A1(\u_cpu.rf_ram.memory[113][2] ),
    .A2(_04388_),
    .ZN(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09659_ (.A1(_04244_),
    .A2(_04384_),
    .B(_04389_),
    .ZN(_00878_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09660_ (.A1(\u_cpu.rf_ram.memory[113][3] ),
    .A2(_04388_),
    .ZN(_04390_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09661_ (.A1(_04247_),
    .A2(_04384_),
    .B(_04390_),
    .ZN(_00879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09662_ (.A1(\u_cpu.rf_ram.memory[113][4] ),
    .A2(_04388_),
    .ZN(_04391_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09663_ (.A1(_04249_),
    .A2(_04384_),
    .B(_04391_),
    .ZN(_00880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09664_ (.A1(\u_cpu.rf_ram.memory[113][5] ),
    .A2(_04388_),
    .ZN(_04392_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09665_ (.A1(_04251_),
    .A2(_04385_),
    .B(_04392_),
    .ZN(_00881_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09666_ (.A1(\u_cpu.rf_ram.memory[113][6] ),
    .A2(_04388_),
    .ZN(_04393_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09667_ (.A1(_04253_),
    .A2(_04385_),
    .B(_04393_),
    .ZN(_00882_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09668_ (.A1(\u_cpu.rf_ram.memory[113][7] ),
    .A2(_04383_),
    .ZN(_04394_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09669_ (.A1(_04255_),
    .A2(_04385_),
    .B(_04394_),
    .ZN(_00883_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09670_ (.I(_03117_),
    .Z(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09671_ (.I(_04395_),
    .Z(_04396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09672_ (.I(_03117_),
    .Z(_04397_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09673_ (.I(_04397_),
    .Z(_04398_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09674_ (.I0(\u_arbiter.i_wb_cpu_rdt[11] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[11] ),
    .S(_01437_),
    .Z(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09675_ (.I0(\u_arbiter.i_wb_cpu_rdt[10] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[10] ),
    .S(_01438_),
    .Z(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09676_ (.I0(\u_arbiter.i_wb_cpu_rdt[9] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ),
    .S(_01437_),
    .Z(_04401_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09677_ (.I0(\u_arbiter.i_wb_cpu_rdt[7] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ),
    .S(_01438_),
    .Z(_04402_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _09678_ (.A1(_04399_),
    .A2(_04400_),
    .A3(_04401_),
    .A4(_04402_),
    .ZN(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09679_ (.I(_03114_),
    .Z(_04404_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09680_ (.I(_01439_),
    .Z(_04405_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09681_ (.A1(_04405_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ),
    .Z(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09682_ (.A1(_04404_),
    .A2(\u_arbiter.i_wb_cpu_rdt[8] ),
    .B(_04406_),
    .ZN(_04407_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09683_ (.A1(_04403_),
    .A2(_04407_),
    .Z(_04408_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09684_ (.I(_04408_),
    .ZN(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09685_ (.A1(_01440_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ),
    .Z(_04410_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09686_ (.A1(_04404_),
    .A2(\u_arbiter.i_wb_cpu_rdt[12] ),
    .B(_04410_),
    .ZN(_04411_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09687_ (.A1(_04409_),
    .A2(_04411_),
    .ZN(_04412_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09688_ (.I(_01437_),
    .Z(_04413_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09689_ (.A1(_04413_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ),
    .Z(_04414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09690_ (.A1(_03114_),
    .A2(\u_arbiter.i_wb_cpu_rdt[0] ),
    .B(_04414_),
    .ZN(_04415_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09691_ (.I(_04415_),
    .Z(_04416_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09692_ (.I(_04413_),
    .Z(_04417_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09693_ (.I0(\u_arbiter.i_wb_cpu_rdt[1] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ),
    .S(_04417_),
    .Z(_04418_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09694_ (.I(_04418_),
    .Z(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09695_ (.I0(\u_arbiter.i_wb_cpu_rdt[6] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ),
    .S(_04417_),
    .Z(_04420_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09696_ (.I(_04420_),
    .ZN(_04421_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09697_ (.A1(_04405_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ),
    .Z(_04422_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09698_ (.A1(_03114_),
    .A2(\u_arbiter.i_wb_cpu_rdt[5] ),
    .B(_04422_),
    .ZN(_04423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09699_ (.A1(_04405_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[3] ),
    .ZN(_04424_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09700_ (.A1(_04405_),
    .A2(_04310_),
    .B(_04424_),
    .ZN(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09701_ (.I0(\u_arbiter.i_wb_cpu_rdt[4] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ),
    .S(_04417_),
    .Z(_04426_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09702_ (.I0(\u_arbiter.i_wb_cpu_rdt[2] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[2] ),
    .S(_04417_),
    .Z(_04427_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09703_ (.A1(_04425_),
    .A2(_04426_),
    .A3(_04427_),
    .ZN(_04428_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09704_ (.A1(_04421_),
    .A2(_04423_),
    .A3(_04428_),
    .ZN(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09705_ (.A1(_04413_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ),
    .Z(_04430_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09706_ (.A1(_03114_),
    .A2(\u_arbiter.i_wb_cpu_rdt[14] ),
    .B(_04430_),
    .ZN(_04431_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09707_ (.I0(\u_arbiter.i_wb_cpu_rdt[15] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ),
    .S(_01439_),
    .Z(_04432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09708_ (.A1(_04431_),
    .A2(_04432_),
    .ZN(_04433_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09709_ (.A1(_04429_),
    .A2(_04433_),
    .ZN(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09710_ (.A1(_04416_),
    .A2(_04419_),
    .A3(_04434_),
    .ZN(_04435_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09711_ (.I(_04427_),
    .Z(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09712_ (.I0(\u_arbiter.i_wb_cpu_rdt[0] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ),
    .S(_01439_),
    .Z(_04437_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09713_ (.A1(_04437_),
    .A2(_04418_),
    .ZN(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09714_ (.I0(\u_arbiter.i_wb_cpu_rdt[14] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ),
    .S(_04413_),
    .Z(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09715_ (.A1(_01438_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ),
    .Z(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09716_ (.A1(_03113_),
    .A2(\u_arbiter.i_wb_cpu_rdt[15] ),
    .B(_04440_),
    .ZN(_04441_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09717_ (.I(_04441_),
    .Z(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09718_ (.A1(_04439_),
    .A2(_04442_),
    .ZN(_04443_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09719_ (.A1(_04437_),
    .A2(_04418_),
    .ZN(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09720_ (.A1(_04443_),
    .A2(_04444_),
    .ZN(_04445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09721_ (.A1(_04438_),
    .A2(_04445_),
    .ZN(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09722_ (.I(_04446_),
    .Z(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09723_ (.A1(_04436_),
    .A2(_04447_),
    .ZN(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09724_ (.A1(_01438_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ),
    .Z(_04449_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09725_ (.A1(_03113_),
    .A2(\u_arbiter.i_wb_cpu_rdt[13] ),
    .B(_04449_),
    .ZN(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09726_ (.A1(_04439_),
    .A2(_04450_),
    .ZN(_04451_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09727_ (.I(_04451_),
    .Z(_04452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09728_ (.A1(_04439_),
    .A2(_04441_),
    .ZN(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09729_ (.I0(\u_arbiter.i_wb_cpu_rdt[8] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ),
    .S(_01439_),
    .Z(_04454_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09730_ (.A1(_04403_),
    .A2(_04454_),
    .Z(_04455_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _09731_ (.A1(_04450_),
    .A2(_04453_),
    .A3(_04455_),
    .ZN(_04456_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09732_ (.I(_04456_),
    .Z(_04457_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09733_ (.A1(_04416_),
    .A2(_04418_),
    .ZN(_04458_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09734_ (.I(_04458_),
    .Z(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09735_ (.A1(_04452_),
    .A2(_04457_),
    .B(_04459_),
    .ZN(_04460_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09736_ (.A1(_04412_),
    .A2(_04435_),
    .B(_04448_),
    .C(_04460_),
    .ZN(_04461_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09737_ (.A1(_04398_),
    .A2(_04461_),
    .ZN(_04462_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09738_ (.A1(_02616_),
    .A2(_04396_),
    .B(_04462_),
    .ZN(_00884_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09739_ (.A1(_04404_),
    .A2(\u_arbiter.i_wb_cpu_ibus_adr[1] ),
    .ZN(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09740_ (.A1(net8),
    .A2(_01433_),
    .A3(_04463_),
    .ZN(_04464_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09741_ (.I(_04464_),
    .Z(_04465_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09742_ (.I(_04465_),
    .Z(_04466_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09743_ (.I(_04466_),
    .Z(_04467_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09744_ (.I(_04425_),
    .Z(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09745_ (.I(_04446_),
    .Z(_04469_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09746_ (.I(_04437_),
    .Z(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09747_ (.A1(_04405_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ),
    .Z(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09748_ (.A1(_04404_),
    .A2(\u_arbiter.i_wb_cpu_rdt[1] ),
    .B(_04471_),
    .ZN(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09749_ (.A1(_04470_),
    .A2(_04472_),
    .ZN(_04473_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09750_ (.I(_04473_),
    .Z(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09751_ (.I(_04431_),
    .Z(_04475_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09752_ (.I0(\u_arbiter.i_wb_cpu_rdt[13] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ),
    .S(_04413_),
    .Z(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09753_ (.I(_04476_),
    .Z(_04477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09754_ (.A1(_04475_),
    .A2(_04477_),
    .ZN(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09755_ (.A1(_04474_),
    .A2(_04478_),
    .ZN(_04479_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09756_ (.A1(_04468_),
    .A2(_04469_),
    .B(_04479_),
    .ZN(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09757_ (.I(_04464_),
    .Z(_04481_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09758_ (.I(_04481_),
    .Z(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09759_ (.A1(_02680_),
    .A2(_04482_),
    .ZN(_04483_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09760_ (.A1(_04467_),
    .A2(_04480_),
    .B(_04483_),
    .ZN(_00885_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09761_ (.I(_04470_),
    .Z(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09762_ (.I(_04475_),
    .Z(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09763_ (.I(_04472_),
    .Z(_04486_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09764_ (.A1(_04429_),
    .A2(_04442_),
    .Z(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _09765_ (.A1(_04412_),
    .A2(_04486_),
    .A3(_04487_),
    .Z(_04488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09766_ (.I(_04439_),
    .Z(_04489_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09767_ (.I(_04432_),
    .Z(_04490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09768_ (.A1(_04489_),
    .A2(_04490_),
    .ZN(_04491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09769_ (.A1(_04478_),
    .A2(_04491_),
    .ZN(_04492_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09770_ (.A1(_04438_),
    .A2(_04445_),
    .Z(_04493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09771_ (.A1(_03118_),
    .A2(_04493_),
    .ZN(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09772_ (.A1(_04484_),
    .A2(_04492_),
    .B(_04494_),
    .ZN(_04495_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09773_ (.A1(_04484_),
    .A2(_04485_),
    .B(_04488_),
    .C(_04495_),
    .ZN(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09774_ (.I(_04426_),
    .Z(_04497_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09775_ (.A1(_04464_),
    .A2(_04493_),
    .ZN(_04498_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09776_ (.I(_04498_),
    .Z(_04499_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09777_ (.I(_04499_),
    .Z(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09778_ (.A1(_02675_),
    .A2(_04482_),
    .B1(_04497_),
    .B2(_04500_),
    .ZN(_04501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09779_ (.A1(_04496_),
    .A2(_04501_),
    .ZN(_00886_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09780_ (.A1(_04433_),
    .A2(_04476_),
    .ZN(_04502_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09781_ (.I(_04502_),
    .Z(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09782_ (.I(_04399_),
    .Z(_04504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09783_ (.I(_04400_),
    .Z(_04505_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09784_ (.A1(_04504_),
    .A2(_04505_),
    .Z(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _09785_ (.A1(_04503_),
    .A2(_04506_),
    .B(_04457_),
    .C(_04492_),
    .ZN(_04507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09786_ (.A1(_04459_),
    .A2(_04507_),
    .ZN(_04508_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09787_ (.I(_04442_),
    .Z(_04509_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09788_ (.I(_04509_),
    .Z(_04510_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09789_ (.I(_04481_),
    .Z(_04511_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09790_ (.A1(_04416_),
    .A2(_04510_),
    .B1(_04447_),
    .B2(_04423_),
    .C(_04511_),
    .ZN(_04512_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09791_ (.A1(_02633_),
    .A2(_04482_),
    .B1(_04508_),
    .B2(_04512_),
    .ZN(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09792_ (.I(_04513_),
    .ZN(_00887_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09793_ (.I(_04421_),
    .Z(_04514_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09794_ (.A1(_02676_),
    .A2(_04395_),
    .ZN(_04515_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09795_ (.A1(_04435_),
    .A2(_04495_),
    .B1(_04500_),
    .B2(_04514_),
    .C(_04515_),
    .ZN(_00888_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09796_ (.I(_03118_),
    .Z(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09797_ (.A1(_04415_),
    .A2(_04418_),
    .ZN(_04517_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09798_ (.I(_04517_),
    .Z(_04518_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09799_ (.A1(_04475_),
    .A2(_04442_),
    .ZN(_04519_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09800_ (.I(_04519_),
    .Z(_04520_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09801_ (.A1(_04514_),
    .A2(_04423_),
    .B(_04506_),
    .ZN(_04521_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09802_ (.A1(_04431_),
    .A2(_04442_),
    .ZN(_04522_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09803_ (.I(_04522_),
    .Z(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _09804_ (.A1(_04436_),
    .A2(_04457_),
    .B1(_04503_),
    .B2(_04521_),
    .C1(_04523_),
    .C2(_04477_),
    .ZN(_04524_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09805_ (.I(_04473_),
    .Z(_04525_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09806_ (.I(_04446_),
    .Z(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09807_ (.I0(\u_arbiter.i_wb_cpu_rdt[12] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ),
    .S(_04417_),
    .Z(_04527_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09808_ (.I(_04527_),
    .Z(_04528_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09809_ (.A1(_04526_),
    .A2(_04479_),
    .B(_04528_),
    .ZN(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _09810_ (.A1(_04518_),
    .A2(_04520_),
    .B1(_04524_),
    .B2(_04525_),
    .C(_04529_),
    .ZN(_04530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09811_ (.A1(_04516_),
    .A2(_04530_),
    .ZN(_04531_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09812_ (.A1(_02557_),
    .A2(_04396_),
    .B(_04531_),
    .ZN(_00889_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09813_ (.A1(_04411_),
    .A2(_04478_),
    .ZN(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09814_ (.A1(_04504_),
    .A2(_04502_),
    .ZN(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09815_ (.A1(_04505_),
    .A2(_04514_),
    .B(_04533_),
    .ZN(_04534_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _09816_ (.A1(_04468_),
    .A2(_04457_),
    .B(_04532_),
    .C(_04534_),
    .ZN(_04535_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _09817_ (.A1(_04484_),
    .A2(_04485_),
    .B1(_04525_),
    .B2(_04535_),
    .C(_04493_),
    .ZN(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09818_ (.A1(_04493_),
    .A2(_04477_),
    .B(_04536_),
    .C(_04395_),
    .ZN(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09819_ (.A1(_02671_),
    .A2(_04396_),
    .B(_04537_),
    .ZN(_00890_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09820_ (.A1(_04421_),
    .A2(_04423_),
    .A3(_04506_),
    .Z(_04538_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09821_ (.I(_04538_),
    .ZN(_04539_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09822_ (.A1(_04497_),
    .A2(_04457_),
    .B1(_04503_),
    .B2(_04539_),
    .C(_04532_),
    .ZN(_04540_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09823_ (.A1(_04485_),
    .A2(_04438_),
    .B1(_04525_),
    .B2(_04540_),
    .ZN(_04541_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09824_ (.A1(_04516_),
    .A2(_04541_),
    .ZN(_04542_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09825_ (.A1(_01409_),
    .A2(_04396_),
    .B(_04542_),
    .ZN(_00891_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09826_ (.I0(\u_arbiter.i_wb_cpu_rdt[20] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[4] ),
    .S(_01442_),
    .Z(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09827_ (.A1(_04412_),
    .A2(_04434_),
    .B1(_04453_),
    .B2(_04427_),
    .C(_04486_),
    .ZN(_04544_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09828_ (.I(_04470_),
    .Z(_04545_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09829_ (.I(_04450_),
    .Z(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09830_ (.A1(_04427_),
    .A2(_04546_),
    .A3(_04491_),
    .ZN(_04547_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09831_ (.I(_04451_),
    .Z(_04548_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09832_ (.I(_04527_),
    .Z(_04549_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09833_ (.A1(_04548_),
    .A2(_04456_),
    .B(_04549_),
    .ZN(_04550_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09834_ (.A1(_04545_),
    .A2(_04547_),
    .A3(_04550_),
    .Z(_04551_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09835_ (.A1(_04416_),
    .A2(_04472_),
    .ZN(_04552_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09836_ (.I(_04552_),
    .Z(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09837_ (.A1(_04436_),
    .A2(_04523_),
    .B(_04553_),
    .ZN(_04554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09838_ (.A1(_03118_),
    .A2(_04438_),
    .ZN(_04555_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _09839_ (.A1(_04544_),
    .A2(_04551_),
    .A3(_04554_),
    .A4(_04555_),
    .ZN(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09840_ (.A1(_04499_),
    .A2(_04543_),
    .B(_04556_),
    .ZN(_04557_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09841_ (.A1(_01382_),
    .A2(_04396_),
    .B(_04557_),
    .ZN(_00892_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09842_ (.I(_04498_),
    .Z(_04558_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09843_ (.I0(\u_arbiter.i_wb_cpu_rdt[21] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[5] ),
    .S(_01447_),
    .Z(_04559_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09844_ (.I(_04444_),
    .Z(_04560_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09845_ (.I(_04522_),
    .Z(_04561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09846_ (.A1(_04425_),
    .A2(_04561_),
    .ZN(_04562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09847_ (.A1(_04527_),
    .A2(_04456_),
    .ZN(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09848_ (.A1(_04545_),
    .A2(_04563_),
    .ZN(_04564_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09849_ (.A1(_04475_),
    .A2(_04490_),
    .ZN(_04565_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09850_ (.I(_04565_),
    .Z(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09851_ (.A1(_04432_),
    .A2(_04477_),
    .ZN(_04567_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09852_ (.A1(_04475_),
    .A2(_04567_),
    .ZN(_04568_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09853_ (.A1(_04470_),
    .A2(_04566_),
    .B1(_04568_),
    .B2(_04419_),
    .ZN(_04569_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09854_ (.A1(_04486_),
    .A2(_04564_),
    .B1(_04569_),
    .B2(_04468_),
    .ZN(_04570_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09855_ (.A1(_04560_),
    .A2(_04562_),
    .B(_04570_),
    .ZN(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09856_ (.I(_04397_),
    .Z(_04572_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09857_ (.A1(_04558_),
    .A2(_04559_),
    .B1(_04571_),
    .B2(_04572_),
    .ZN(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09858_ (.A1(_02571_),
    .A2(_04398_),
    .B(_04573_),
    .ZN(_00893_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09859_ (.I0(\u_arbiter.i_wb_cpu_rdt[22] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[6] ),
    .S(_01446_),
    .Z(_04574_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09860_ (.I(_04552_),
    .Z(_04575_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09861_ (.A1(_04525_),
    .A2(_04563_),
    .ZN(_04576_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09862_ (.A1(_04563_),
    .A2(_04568_),
    .ZN(_04577_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09863_ (.A1(_04458_),
    .A2(_04577_),
    .ZN(_04578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09864_ (.A1(_04518_),
    .A2(_04578_),
    .ZN(_04579_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09865_ (.A1(_04497_),
    .A2(_04576_),
    .B(_04579_),
    .ZN(_04580_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09866_ (.A1(_04426_),
    .A2(_04561_),
    .ZN(_04581_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09867_ (.I(_04552_),
    .Z(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09868_ (.A1(_04420_),
    .A2(_04509_),
    .B1(_04443_),
    .B2(_04574_),
    .C(_04582_),
    .ZN(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09869_ (.A1(_04575_),
    .A2(_04580_),
    .B1(_04581_),
    .B2(_04583_),
    .ZN(_04584_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09870_ (.A1(_04481_),
    .A2(_04526_),
    .ZN(_04585_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09871_ (.A1(_04558_),
    .A2(_04574_),
    .B1(_04584_),
    .B2(_04585_),
    .ZN(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09872_ (.A1(_02562_),
    .A2(_04398_),
    .B(_04586_),
    .ZN(_00894_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09873_ (.A1(_02722_),
    .A2(_04224_),
    .ZN(_04587_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09874_ (.I(_04587_),
    .Z(_04588_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09875_ (.I(_04587_),
    .Z(_04589_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09876_ (.A1(\u_cpu.rf_ram.memory[114][0] ),
    .A2(_04589_),
    .ZN(_04590_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09877_ (.A1(_04237_),
    .A2(_04588_),
    .B(_04590_),
    .ZN(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09878_ (.A1(\u_cpu.rf_ram.memory[114][1] ),
    .A2(_04589_),
    .ZN(_04591_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09879_ (.A1(_04242_),
    .A2(_04588_),
    .B(_04591_),
    .ZN(_00896_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09880_ (.I(_04587_),
    .Z(_04592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09881_ (.A1(\u_cpu.rf_ram.memory[114][2] ),
    .A2(_04592_),
    .ZN(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09882_ (.A1(_04244_),
    .A2(_04588_),
    .B(_04593_),
    .ZN(_00897_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09883_ (.A1(\u_cpu.rf_ram.memory[114][3] ),
    .A2(_04592_),
    .ZN(_04594_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09884_ (.A1(_04247_),
    .A2(_04588_),
    .B(_04594_),
    .ZN(_00898_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09885_ (.A1(\u_cpu.rf_ram.memory[114][4] ),
    .A2(_04592_),
    .ZN(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09886_ (.A1(_04249_),
    .A2(_04588_),
    .B(_04595_),
    .ZN(_00899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09887_ (.A1(\u_cpu.rf_ram.memory[114][5] ),
    .A2(_04592_),
    .ZN(_04596_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09888_ (.A1(_04251_),
    .A2(_04589_),
    .B(_04596_),
    .ZN(_00900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09889_ (.A1(\u_cpu.rf_ram.memory[114][6] ),
    .A2(_04592_),
    .ZN(_04597_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09890_ (.A1(_04253_),
    .A2(_04589_),
    .B(_04597_),
    .ZN(_00901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09891_ (.A1(\u_cpu.rf_ram.memory[114][7] ),
    .A2(_04587_),
    .ZN(_04598_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09892_ (.A1(_04255_),
    .A2(_04589_),
    .B(_04598_),
    .ZN(_00902_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09893_ (.I0(\u_arbiter.i_wb_cpu_rdt[26] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[10] ),
    .S(_01441_),
    .Z(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09894_ (.A1(_04499_),
    .A2(_04599_),
    .ZN(_04600_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09895_ (.I0(\u_arbiter.i_wb_cpu_rdt[5] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ),
    .S(_01440_),
    .Z(_04601_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09896_ (.I(_04454_),
    .Z(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09897_ (.A1(_04403_),
    .A2(_04602_),
    .ZN(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09898_ (.A1(_04546_),
    .A2(_04453_),
    .ZN(_04604_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09899_ (.A1(_04549_),
    .A2(_04455_),
    .B(_04604_),
    .ZN(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09900_ (.I(_04605_),
    .ZN(_04606_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09901_ (.A1(_04601_),
    .A2(_04603_),
    .B(_04606_),
    .ZN(_04607_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09902_ (.I(_04402_),
    .Z(_04608_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09903_ (.A1(_04489_),
    .A2(_04432_),
    .ZN(_04609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09904_ (.A1(_04546_),
    .A2(_04609_),
    .ZN(_04610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09905_ (.A1(_04527_),
    .A2(_04489_),
    .ZN(_04611_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09906_ (.I(_04611_),
    .ZN(_04612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09907_ (.A1(_04443_),
    .A2(_04546_),
    .ZN(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09908_ (.A1(_04399_),
    .A2(_04527_),
    .ZN(_04614_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09909_ (.A1(_04400_),
    .A2(_04613_),
    .A3(_04614_),
    .ZN(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09910_ (.A1(_04567_),
    .A2(_04612_),
    .B(_04615_),
    .ZN(_04616_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09911_ (.A1(_04610_),
    .A2(_04616_),
    .ZN(_04617_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09912_ (.A1(_04608_),
    .A2(_04548_),
    .B1(_04561_),
    .B2(_04601_),
    .C(_04617_),
    .ZN(_04618_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09913_ (.A1(_04528_),
    .A2(_04610_),
    .B(_04459_),
    .ZN(_04619_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09914_ (.A1(_04607_),
    .A2(_04618_),
    .B(_04619_),
    .ZN(_04620_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09915_ (.A1(_04436_),
    .A2(_04566_),
    .B1(_04523_),
    .B2(_04608_),
    .C(_04472_),
    .ZN(_04621_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09916_ (.A1(_04484_),
    .A2(_04621_),
    .ZN(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _09917_ (.A1(_04485_),
    .A2(_04601_),
    .B1(_04433_),
    .B2(_04599_),
    .C1(_04520_),
    .C2(_04608_),
    .ZN(_04623_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09918_ (.A1(_04444_),
    .A2(_04623_),
    .ZN(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09919_ (.A1(_04620_),
    .A2(_04622_),
    .B(_04624_),
    .C(_04585_),
    .ZN(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09920_ (.A1(_04600_),
    .A2(_04625_),
    .Z(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09921_ (.A1(_01381_),
    .A2(_04398_),
    .B(_04626_),
    .ZN(_00903_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09922_ (.A1(_02679_),
    .A2(_02703_),
    .A3(_01377_),
    .B(_02529_),
    .ZN(_04627_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09923_ (.A1(_04465_),
    .A2(_04627_),
    .Z(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09924_ (.I(_04628_),
    .Z(_04629_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09925_ (.I(_04481_),
    .Z(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09926_ (.A1(\u_cpu.cpu.immdec.imm24_20[1] ),
    .A2(_04630_),
    .ZN(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09927_ (.A1(\u_cpu.cpu.immdec.imm24_20[0] ),
    .A2(_04628_),
    .ZN(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09928_ (.A1(_04629_),
    .A2(_04631_),
    .B(_04632_),
    .C(_04557_),
    .ZN(_00904_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09929_ (.A1(_04397_),
    .A2(_04627_),
    .ZN(_04633_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09930_ (.A1(\u_cpu.cpu.immdec.imm24_20[1] ),
    .A2(_04629_),
    .B1(_04633_),
    .B2(\u_cpu.cpu.immdec.imm24_20[2] ),
    .ZN(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09931_ (.A1(_04573_),
    .A2(_04634_),
    .ZN(_00905_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09932_ (.I(\u_cpu.cpu.immdec.imm24_20[2] ),
    .ZN(_04635_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09933_ (.I(_04481_),
    .Z(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09934_ (.A1(\u_cpu.cpu.immdec.imm24_20[3] ),
    .A2(_04627_),
    .B(_04636_),
    .ZN(_04637_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09935_ (.A1(_04635_),
    .A2(_04629_),
    .B1(_04637_),
    .B2(_04586_),
    .ZN(_00906_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09936_ (.I0(\u_arbiter.i_wb_cpu_rdt[23] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[7] ),
    .S(_01441_),
    .Z(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09937_ (.A1(_04549_),
    .A2(_04456_),
    .B1(_04502_),
    .B2(_04506_),
    .ZN(_04639_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09938_ (.A1(_04578_),
    .A2(_04639_),
    .B(_04423_),
    .ZN(_04640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09939_ (.A1(_04579_),
    .A2(_04640_),
    .ZN(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09940_ (.I(_04489_),
    .Z(_04642_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09941_ (.A1(_04505_),
    .A2(_04490_),
    .Z(_04643_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09942_ (.A1(_04642_),
    .A2(_04638_),
    .B(_04643_),
    .C(_04520_),
    .ZN(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09943_ (.A1(_04601_),
    .A2(_04609_),
    .B(_04553_),
    .ZN(_04645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09944_ (.A1(_04582_),
    .A2(_04641_),
    .B1(_04644_),
    .B2(_04645_),
    .C(_04526_),
    .ZN(_04646_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09945_ (.A1(_04469_),
    .A2(_04638_),
    .B(_04646_),
    .C(_04466_),
    .ZN(_04647_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09946_ (.A1(\u_cpu.cpu.immdec.imm24_20[4] ),
    .A2(_04572_),
    .ZN(_04648_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09947_ (.A1(\u_cpu.cpu.immdec.imm24_20[3] ),
    .A2(_04629_),
    .ZN(_04649_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09948_ (.A1(_04629_),
    .A2(_04647_),
    .A3(_04648_),
    .B(_04649_),
    .ZN(_00907_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09949_ (.I(_04504_),
    .Z(_04650_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09950_ (.A1(_04650_),
    .A2(_04452_),
    .B1(_04507_),
    .B2(_04420_),
    .C(_04564_),
    .ZN(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09951_ (.I(_04443_),
    .Z(_04652_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09952_ (.I0(\u_arbiter.i_wb_cpu_rdt[24] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[8] ),
    .S(_01446_),
    .Z(_04653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09953_ (.A1(_04650_),
    .A2(_04510_),
    .B1(_04652_),
    .B2(_04653_),
    .ZN(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09954_ (.A1(_04419_),
    .A2(_04514_),
    .B1(_04560_),
    .B2(_04654_),
    .ZN(_04655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09955_ (.A1(_04585_),
    .A2(_04655_),
    .ZN(_04656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _09956_ (.A1(\u_cpu.cpu.immdec.imm24_20[4] ),
    .A2(_04628_),
    .B1(_04633_),
    .B2(\u_cpu.cpu.immdec.imm30_25[0] ),
    .C1(_04653_),
    .C2(_04558_),
    .ZN(_04657_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09957_ (.A1(_04651_),
    .A2(_04656_),
    .B(_04657_),
    .ZN(_00908_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09958_ (.A1(_04470_),
    .A2(_04485_),
    .ZN(_04658_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09959_ (.A1(_04546_),
    .A2(_04603_),
    .ZN(_04659_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09960_ (.A1(_04492_),
    .A2(_04659_),
    .B(_04427_),
    .ZN(_04660_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09961_ (.A1(_04528_),
    .A2(_04567_),
    .B(_04615_),
    .ZN(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09962_ (.A1(_04545_),
    .A2(_04563_),
    .A3(_04660_),
    .A4(_04661_),
    .ZN(_04662_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _09963_ (.A1(_04528_),
    .A2(_04484_),
    .B1(_04486_),
    .B2(_04658_),
    .C(_04662_),
    .ZN(_04663_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09964_ (.A1(_04585_),
    .A2(_04663_),
    .Z(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09965_ (.A1(_02679_),
    .A2(_02703_),
    .A3(_02677_),
    .ZN(_04665_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09966_ (.A1(_02529_),
    .A2(_04665_),
    .ZN(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09967_ (.A1(_04465_),
    .A2(_04666_),
    .ZN(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09968_ (.A1(_03115_),
    .A2(\u_arbiter.i_wb_cpu_rdt[25] ),
    .ZN(_04668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09969_ (.A1(_01443_),
    .A2(\u_arbiter.i_wb_cpu_rdt[9] ),
    .ZN(_04669_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09970_ (.A1(_04498_),
    .A2(_04668_),
    .A3(_04669_),
    .ZN(_04670_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09971_ (.A1(\u_cpu.cpu.immdec.imm30_25[1] ),
    .A2(_04516_),
    .B(_04667_),
    .C(_04670_),
    .ZN(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09972_ (.A1(_04465_),
    .A2(_04666_),
    .Z(_04672_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09973_ (.A1(\u_cpu.cpu.immdec.imm30_25[0] ),
    .A2(_04672_),
    .ZN(_04673_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09974_ (.A1(_04664_),
    .A2(_04671_),
    .B(_04673_),
    .ZN(_00909_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09975_ (.A1(_04397_),
    .A2(_04666_),
    .ZN(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09976_ (.A1(\u_cpu.cpu.immdec.imm30_25[1] ),
    .A2(_04672_),
    .B1(_04674_),
    .B2(\u_cpu.cpu.immdec.imm30_25[2] ),
    .ZN(_04675_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09977_ (.A1(_04626_),
    .A2(_04675_),
    .ZN(_00910_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09978_ (.A1(_04563_),
    .A2(_04661_),
    .ZN(_04676_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09979_ (.A1(_04425_),
    .A2(_04566_),
    .A3(_04659_),
    .ZN(_04677_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09980_ (.A1(_04545_),
    .A2(_04677_),
    .ZN(_04678_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09981_ (.A1(_04420_),
    .A2(_04492_),
    .B(_04676_),
    .C(_04678_),
    .ZN(_04679_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09982_ (.I(_04602_),
    .Z(_04680_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09983_ (.A1(_04468_),
    .A2(_04566_),
    .B1(_04523_),
    .B2(_04680_),
    .C(_04486_),
    .ZN(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09984_ (.I0(\u_arbiter.i_wb_cpu_rdt[27] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[11] ),
    .S(_01446_),
    .Z(_04682_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09985_ (.A1(_04680_),
    .A2(_04609_),
    .B1(_04682_),
    .B2(_04652_),
    .C(_04575_),
    .ZN(_04683_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _09986_ (.A1(_04494_),
    .A2(_04679_),
    .A3(_04681_),
    .A4(_04683_),
    .Z(_04684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _09987_ (.A1(\u_cpu.cpu.immdec.imm30_25[2] ),
    .A2(_04672_),
    .B1(_04674_),
    .B2(\u_cpu.cpu.immdec.imm30_25[3] ),
    .C1(_04682_),
    .C2(_04558_),
    .ZN(_04685_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09988_ (.A1(_04684_),
    .A2(_04685_),
    .ZN(_00911_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09989_ (.A1(_01443_),
    .A2(\u_arbiter.i_wb_cpu_rdt[12] ),
    .Z(_04686_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09990_ (.A1(_03115_),
    .A2(\u_arbiter.i_wb_cpu_rdt[28] ),
    .B(_04686_),
    .ZN(_04687_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09991_ (.A1(_04497_),
    .A2(_04603_),
    .B(_04606_),
    .ZN(_04688_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09992_ (.A1(_04401_),
    .A2(_04452_),
    .B1(_04523_),
    .B2(_04528_),
    .C(_04617_),
    .ZN(_04689_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09993_ (.A1(_04688_),
    .A2(_04689_),
    .B(_04619_),
    .ZN(_04690_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09994_ (.A1(_01440_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ),
    .Z(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09995_ (.A1(_03115_),
    .A2(\u_arbiter.i_wb_cpu_rdt[9] ),
    .B(_04691_),
    .ZN(_04692_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09996_ (.A1(_04692_),
    .A2(_04575_),
    .A3(_04520_),
    .ZN(_04693_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09997_ (.A1(_04494_),
    .A2(_04690_),
    .A3(_04693_),
    .ZN(_04694_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09998_ (.A1(_02530_),
    .A2(_04465_),
    .A3(_04665_),
    .ZN(_04695_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09999_ (.A1(\u_cpu.cpu.immdec.imm30_25[3] ),
    .A2(_04667_),
    .B1(_04695_),
    .B2(\u_cpu.cpu.immdec.imm30_25[4] ),
    .ZN(_04696_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10000_ (.A1(_04500_),
    .A2(_04687_),
    .B(_04694_),
    .C(_04696_),
    .ZN(_00912_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10001_ (.A1(_01443_),
    .A2(\u_arbiter.i_wb_cpu_rdt[13] ),
    .Z(_04697_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10002_ (.A1(_03115_),
    .A2(\u_arbiter.i_wb_cpu_rdt[29] ),
    .B(_04697_),
    .ZN(_04698_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10003_ (.A1(_04642_),
    .A2(_04582_),
    .ZN(_04699_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10004_ (.I(_04610_),
    .Z(_04700_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10005_ (.I(_04505_),
    .Z(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10006_ (.A1(_04701_),
    .A2(_04548_),
    .B(_04615_),
    .C(_04612_),
    .ZN(_04702_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10007_ (.A1(_04700_),
    .A2(_04702_),
    .B(_04619_),
    .ZN(_04703_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10008_ (.A1(_04643_),
    .A2(_04699_),
    .B(_04703_),
    .C(_04555_),
    .ZN(_04704_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10009_ (.A1(\u_cpu.cpu.immdec.imm30_25[4] ),
    .A2(_04667_),
    .B1(_04695_),
    .B2(\u_cpu.cpu.immdec.imm30_25[5] ),
    .ZN(_04705_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10010_ (.A1(_04500_),
    .A2(_04698_),
    .B(_04704_),
    .C(_04705_),
    .ZN(_00913_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10011_ (.I0(\u_arbiter.i_wb_cpu_rdt[30] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[14] ),
    .S(_01447_),
    .Z(_04706_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10012_ (.A1(_04505_),
    .A2(_04411_),
    .B(_04504_),
    .ZN(_04707_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _10013_ (.A1(_04504_),
    .A2(_04701_),
    .B1(_04538_),
    .B2(_04707_),
    .C(_04503_),
    .ZN(_04708_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10014_ (.A1(_04477_),
    .A2(_04519_),
    .ZN(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10015_ (.I(_04709_),
    .Z(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10016_ (.A1(_04680_),
    .A2(_04452_),
    .B(_04710_),
    .C(_04612_),
    .ZN(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10017_ (.A1(_04708_),
    .A2(_04711_),
    .B(_04619_),
    .ZN(_04712_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10018_ (.A1(_04499_),
    .A2(_04706_),
    .B1(_04712_),
    .B2(_04395_),
    .ZN(_04713_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10019_ (.A1(\u_cpu.cpu.immdec.imm30_25[5] ),
    .A2(_04672_),
    .ZN(_04714_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10020_ (.I(\u_cpu.cpu.immdec.imm19_12_20[0] ),
    .ZN(_04715_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10021_ (.A1(_02675_),
    .A2(_02703_),
    .B(_02680_),
    .ZN(_04716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10022_ (.A1(_02625_),
    .A2(_04716_),
    .ZN(_04717_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10023_ (.A1(_04715_),
    .A2(_04716_),
    .B(_04717_),
    .C(_02682_),
    .ZN(_04718_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10024_ (.A1(\u_cpu.cpu.immdec.imm7 ),
    .A2(_02682_),
    .B(_04674_),
    .C(_04718_),
    .ZN(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10025_ (.A1(_04713_),
    .A2(_04714_),
    .A3(_04719_),
    .ZN(_00914_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10026_ (.A1(_01440_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ),
    .Z(_04720_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10027_ (.A1(_04404_),
    .A2(\u_arbiter.i_wb_cpu_rdt[7] ),
    .B(_04720_),
    .ZN(_04721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10028_ (.A1(_04487_),
    .A2(_04491_),
    .ZN(_04722_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10029_ (.A1(_04409_),
    .A2(_04549_),
    .A3(_04434_),
    .ZN(_04723_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10030_ (.A1(_04721_),
    .A2(_04722_),
    .B(_04723_),
    .C(_04419_),
    .ZN(_04724_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10031_ (.A1(_04549_),
    .A2(_04561_),
    .ZN(_04725_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10032_ (.A1(_04721_),
    .A2(_04489_),
    .ZN(_04726_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10033_ (.A1(_04402_),
    .A2(_04502_),
    .B1(_04726_),
    .B2(_04509_),
    .ZN(_04727_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10034_ (.A1(_04721_),
    .A2(_04710_),
    .B1(_04725_),
    .B2(_04727_),
    .C(_04474_),
    .ZN(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10035_ (.A1(_04416_),
    .A2(_04724_),
    .B(_04728_),
    .ZN(_04729_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10036_ (.A1(_04436_),
    .A2(_04510_),
    .B1(_04652_),
    .B2(_04608_),
    .C(_04582_),
    .ZN(_04730_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10037_ (.A1(_04729_),
    .A2(_04730_),
    .ZN(_04731_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10038_ (.A1(_04608_),
    .A2(_04499_),
    .B1(_04731_),
    .B2(_04585_),
    .ZN(_04732_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10039_ (.A1(_02674_),
    .A2(_02625_),
    .B(_04466_),
    .ZN(_04733_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10040_ (.A1(\u_cpu.cpu.immdec.imm7 ),
    .A2(_02530_),
    .ZN(_04734_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10041_ (.A1(_04732_),
    .A2(_04733_),
    .B1(_04734_),
    .B2(_04467_),
    .ZN(_00915_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10042_ (.A1(_02605_),
    .A2(_02680_),
    .ZN(_04735_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10043_ (.A1(_02539_),
    .A2(_02624_),
    .A3(_04735_),
    .ZN(_04736_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10044_ (.A1(_02529_),
    .A2(_04736_),
    .B(_03117_),
    .ZN(_04737_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10045_ (.I(_04737_),
    .Z(_04738_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10046_ (.I(_04737_),
    .Z(_04739_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10047_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[1] ),
    .A2(_04636_),
    .B(_04739_),
    .ZN(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10048_ (.A1(_04715_),
    .A2(_04738_),
    .B1(_04740_),
    .B2(_04557_),
    .ZN(_00916_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10049_ (.I(\u_cpu.cpu.immdec.imm19_12_20[1] ),
    .ZN(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10050_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[2] ),
    .A2(_04636_),
    .B(_04737_),
    .ZN(_04742_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10051_ (.A1(_04741_),
    .A2(_04738_),
    .B1(_04742_),
    .B2(_04531_),
    .ZN(_00917_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10052_ (.I(\u_cpu.cpu.immdec.imm19_12_20[2] ),
    .ZN(_04743_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10053_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[3] ),
    .A2(_04636_),
    .B(_04737_),
    .ZN(_04744_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10054_ (.A1(_04743_),
    .A2(_04738_),
    .B1(_04744_),
    .B2(_04537_),
    .ZN(_00918_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10055_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[3] ),
    .A2(_04739_),
    .ZN(_04745_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10056_ (.A1(\u_cpu.cpu.csr_imm ),
    .A2(_02530_),
    .A3(_04482_),
    .A4(_04736_),
    .ZN(_04746_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10057_ (.A1(_04542_),
    .A2(_04745_),
    .A3(_04746_),
    .ZN(_00919_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10058_ (.A1(_04692_),
    .A2(_04709_),
    .B(_04474_),
    .ZN(_04747_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10059_ (.A1(_04509_),
    .A2(_04548_),
    .ZN(_04748_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10060_ (.A1(_04411_),
    .A2(_04429_),
    .A3(_04490_),
    .Z(_04749_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10061_ (.A1(_04517_),
    .A2(_04642_),
    .A3(_04749_),
    .ZN(_04750_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10062_ (.A1(_04747_),
    .A2(_04748_),
    .B(_04750_),
    .ZN(_04751_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10063_ (.A1(_04553_),
    .A2(_04609_),
    .ZN(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10064_ (.A1(_04532_),
    .A2(_04709_),
    .ZN(_04753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10065_ (.A1(_04601_),
    .A2(_04456_),
    .ZN(_04754_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10066_ (.A1(_04721_),
    .A2(_04710_),
    .B1(_04753_),
    .B2(_04754_),
    .C(_04474_),
    .ZN(_04755_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10067_ (.A1(_04752_),
    .A2(_04726_),
    .B(_04755_),
    .C(_04526_),
    .ZN(_04756_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10068_ (.A1(_04721_),
    .A2(_04751_),
    .B(_04756_),
    .ZN(_04757_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10069_ (.A1(_04490_),
    .A2(_04438_),
    .B(_04757_),
    .C(_04572_),
    .ZN(_04758_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10070_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[5] ),
    .A2(_04630_),
    .B(_04739_),
    .ZN(_04759_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10071_ (.A1(_01391_),
    .A2(_04738_),
    .B1(_04758_),
    .B2(_04759_),
    .ZN(_00920_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10072_ (.I0(\u_arbiter.i_wb_cpu_rdt[16] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[0] ),
    .S(_01446_),
    .Z(_04760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10073_ (.A1(_04652_),
    .A2(_04760_),
    .ZN(_04761_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10074_ (.A1(_04602_),
    .A2(_04642_),
    .B(_04553_),
    .C(_04609_),
    .ZN(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10075_ (.A1(_04407_),
    .A2(_04709_),
    .B(_04474_),
    .ZN(_04763_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10076_ (.A1(_04420_),
    .A2(_04455_),
    .B(_04604_),
    .ZN(_04764_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10077_ (.A1(_04561_),
    .A2(_04502_),
    .B(_04602_),
    .ZN(_04765_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10078_ (.A1(_04753_),
    .A2(_04764_),
    .A3(_04765_),
    .ZN(_04766_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10079_ (.A1(_04407_),
    .A2(_04518_),
    .A3(_04749_),
    .B(_04552_),
    .ZN(_04767_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10080_ (.A1(_04763_),
    .A2(_04766_),
    .B(_04767_),
    .C(_04658_),
    .ZN(_04768_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10081_ (.A1(_04761_),
    .A2(_04762_),
    .B(_04447_),
    .C(_04768_),
    .ZN(_04769_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10082_ (.A1(_04469_),
    .A2(_04760_),
    .B(_04769_),
    .C(_04466_),
    .ZN(_04770_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10083_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[6] ),
    .A2(_04572_),
    .ZN(_04771_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10084_ (.I(_04737_),
    .Z(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10085_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[5] ),
    .A2(_04772_),
    .ZN(_04773_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10086_ (.A1(_04738_),
    .A2(_04770_),
    .A3(_04771_),
    .B(_04773_),
    .ZN(_00921_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10087_ (.I0(\u_arbiter.i_wb_cpu_rdt[17] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[1] ),
    .S(_01441_),
    .Z(_04774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10088_ (.A1(_04401_),
    .A2(_04642_),
    .B1(_04443_),
    .B2(_04774_),
    .C(_04553_),
    .ZN(_04775_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10089_ (.A1(_04447_),
    .A2(_04775_),
    .ZN(_04776_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10090_ (.A1(_04550_),
    .A2(_04700_),
    .ZN(_04777_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10091_ (.A1(_04747_),
    .A2(_04777_),
    .ZN(_04778_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10092_ (.A1(_04692_),
    .A2(_04751_),
    .B(_04778_),
    .C(_04575_),
    .ZN(_04779_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10093_ (.A1(_04447_),
    .A2(_04774_),
    .B1(_04776_),
    .B2(_04779_),
    .C(_04511_),
    .ZN(_04780_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10094_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[7] ),
    .A2(_04572_),
    .ZN(_04781_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10095_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[6] ),
    .A2(_04772_),
    .ZN(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10096_ (.A1(_04772_),
    .A2(_04780_),
    .A3(_04781_),
    .B(_04782_),
    .ZN(_00922_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10097_ (.I0(\u_arbiter.i_wb_cpu_rdt[18] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[2] ),
    .S(_01442_),
    .Z(_04783_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10098_ (.A1(_04701_),
    .A2(_04750_),
    .B(_04444_),
    .ZN(_04784_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10099_ (.A1(_04548_),
    .A2(_04565_),
    .B(_04550_),
    .ZN(_04785_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10100_ (.A1(_04701_),
    .A2(_04700_),
    .B(_04785_),
    .C(_04459_),
    .ZN(_04786_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10101_ (.A1(_04784_),
    .A2(_04786_),
    .B(_04699_),
    .ZN(_04787_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10102_ (.A1(_04469_),
    .A2(_04783_),
    .B(_04787_),
    .C(_04511_),
    .ZN(_04788_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10103_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[8] ),
    .A2(_04395_),
    .ZN(_04789_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10104_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[7] ),
    .A2(_04739_),
    .ZN(_04790_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10105_ (.A1(_04772_),
    .A2(_04788_),
    .A3(_04789_),
    .B(_04790_),
    .ZN(_00923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10106_ (.A1(_04650_),
    .A2(_04710_),
    .ZN(_04791_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10107_ (.A1(_04550_),
    .A2(_04791_),
    .ZN(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10108_ (.A1(_01442_),
    .A2(_04310_),
    .ZN(_04793_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10109_ (.A1(_01442_),
    .A2(\u_arbiter.i_wb_cpu_rdt[19] ),
    .B(_04526_),
    .C(_04793_),
    .ZN(_04794_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10110_ (.A1(_04397_),
    .A2(_04794_),
    .ZN(_04795_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10111_ (.A1(_04650_),
    .A2(_04750_),
    .B1(_04792_),
    .B2(_04459_),
    .C(_04795_),
    .ZN(_04796_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10112_ (.A1(_02684_),
    .A2(\u_cpu.cpu.immdec.imm24_20[0] ),
    .ZN(_04797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10113_ (.A1(_04511_),
    .A2(_04797_),
    .ZN(_04798_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10114_ (.A1(_02676_),
    .A2(_02625_),
    .B(_04798_),
    .ZN(_04799_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10115_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[8] ),
    .A2(_04739_),
    .ZN(_04800_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10116_ (.A1(_04772_),
    .A2(_04796_),
    .A3(_04799_),
    .B(_04800_),
    .ZN(_00924_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _10117_ (.A1(_04532_),
    .A2(_04710_),
    .A3(_04615_),
    .A4(_04612_),
    .ZN(_04801_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10118_ (.I0(\u_arbiter.i_wb_cpu_rdt[31] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[15] ),
    .S(_01447_),
    .Z(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10119_ (.A1(\u_cpu.cpu.immdec.imm31 ),
    .A2(_04630_),
    .B1(_04558_),
    .B2(_04802_),
    .ZN(_04803_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10120_ (.A1(_04467_),
    .A2(_04619_),
    .A3(_04801_),
    .B(_04803_),
    .ZN(_00925_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10121_ (.I(\u_cpu.cpu.genblk3.csr.timer_irq_r ),
    .ZN(_04804_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10122_ (.A1(_04026_),
    .A2(_02705_),
    .Z(_04805_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10123_ (.A1(\u_cpu.cpu.genblk3.csr.mie_mtie ),
    .A2(\u_cpu.cpu.genblk3.csr.mstatus_mie ),
    .A3(\u_cpu.cpu.genblk3.csr.i_mtip ),
    .A4(_04805_),
    .ZN(_04806_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10124_ (.A1(_04804_),
    .A2(_04805_),
    .B(_04806_),
    .ZN(_00926_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10125_ (.I(_02738_),
    .Z(_04807_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10126_ (.I(_04807_),
    .Z(_04808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10127_ (.A1(_02890_),
    .A2(_02965_),
    .ZN(_04809_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10128_ (.I(_04809_),
    .Z(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10129_ (.I(_04809_),
    .Z(_04811_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10130_ (.A1(\u_cpu.rf_ram.memory[32][0] ),
    .A2(_04811_),
    .ZN(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10131_ (.A1(_04808_),
    .A2(_04810_),
    .B(_04812_),
    .ZN(_00927_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10132_ (.I(_02744_),
    .Z(_04813_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10133_ (.I(_04813_),
    .Z(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10134_ (.A1(\u_cpu.rf_ram.memory[32][1] ),
    .A2(_04811_),
    .ZN(_04815_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10135_ (.A1(_04814_),
    .A2(_04810_),
    .B(_04815_),
    .ZN(_00928_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10136_ (.I(_02750_),
    .Z(_04816_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10137_ (.I(_04816_),
    .Z(_04817_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10138_ (.I(_04809_),
    .Z(_04818_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10139_ (.A1(\u_cpu.rf_ram.memory[32][2] ),
    .A2(_04818_),
    .ZN(_04819_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10140_ (.A1(_04817_),
    .A2(_04810_),
    .B(_04819_),
    .ZN(_00929_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10141_ (.I(_02756_),
    .Z(_04820_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10142_ (.I(_04820_),
    .Z(_04821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10143_ (.A1(\u_cpu.rf_ram.memory[32][3] ),
    .A2(_04818_),
    .ZN(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10144_ (.A1(_04821_),
    .A2(_04810_),
    .B(_04822_),
    .ZN(_00930_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10145_ (.I(_02761_),
    .Z(_04823_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10146_ (.I(_04823_),
    .Z(_04824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10147_ (.A1(\u_cpu.rf_ram.memory[32][4] ),
    .A2(_04818_),
    .ZN(_04825_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10148_ (.A1(_04824_),
    .A2(_04810_),
    .B(_04825_),
    .ZN(_00931_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10149_ (.I(_02766_),
    .Z(_04826_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10150_ (.I(_04826_),
    .Z(_04827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10151_ (.A1(\u_cpu.rf_ram.memory[32][5] ),
    .A2(_04818_),
    .ZN(_04828_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10152_ (.A1(_04827_),
    .A2(_04811_),
    .B(_04828_),
    .ZN(_00932_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10153_ (.I(_02771_),
    .Z(_04829_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10154_ (.I(_04829_),
    .Z(_04830_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10155_ (.A1(\u_cpu.rf_ram.memory[32][6] ),
    .A2(_04818_),
    .ZN(_04831_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10156_ (.A1(_04830_),
    .A2(_04811_),
    .B(_04831_),
    .ZN(_00933_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10157_ (.I(_02776_),
    .Z(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10158_ (.I(_04832_),
    .Z(_04833_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10159_ (.A1(\u_cpu.rf_ram.memory[32][7] ),
    .A2(_04809_),
    .ZN(_04834_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10160_ (.A1(_04833_),
    .A2(_04811_),
    .B(_04834_),
    .ZN(_00934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10161_ (.A1(_03367_),
    .A2(_03062_),
    .ZN(_04835_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10162_ (.I(_04835_),
    .Z(_04836_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10163_ (.I(_04835_),
    .Z(_04837_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10164_ (.A1(\u_cpu.rf_ram.memory[31][0] ),
    .A2(_04837_),
    .ZN(_04838_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10165_ (.A1(_04808_),
    .A2(_04836_),
    .B(_04838_),
    .ZN(_00935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10166_ (.A1(\u_cpu.rf_ram.memory[31][1] ),
    .A2(_04837_),
    .ZN(_04839_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10167_ (.A1(_04814_),
    .A2(_04836_),
    .B(_04839_),
    .ZN(_00936_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10168_ (.I(_04835_),
    .Z(_04840_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10169_ (.A1(\u_cpu.rf_ram.memory[31][2] ),
    .A2(_04840_),
    .ZN(_04841_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10170_ (.A1(_04817_),
    .A2(_04836_),
    .B(_04841_),
    .ZN(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10171_ (.A1(\u_cpu.rf_ram.memory[31][3] ),
    .A2(_04840_),
    .ZN(_04842_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10172_ (.A1(_04821_),
    .A2(_04836_),
    .B(_04842_),
    .ZN(_00938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10173_ (.A1(\u_cpu.rf_ram.memory[31][4] ),
    .A2(_04840_),
    .ZN(_04843_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10174_ (.A1(_04824_),
    .A2(_04836_),
    .B(_04843_),
    .ZN(_00939_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10175_ (.A1(\u_cpu.rf_ram.memory[31][5] ),
    .A2(_04840_),
    .ZN(_04844_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10176_ (.A1(_04827_),
    .A2(_04837_),
    .B(_04844_),
    .ZN(_00940_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10177_ (.A1(\u_cpu.rf_ram.memory[31][6] ),
    .A2(_04840_),
    .ZN(_04845_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10178_ (.A1(_04830_),
    .A2(_04837_),
    .B(_04845_),
    .ZN(_00941_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10179_ (.A1(\u_cpu.rf_ram.memory[31][7] ),
    .A2(_04835_),
    .ZN(_04846_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10180_ (.A1(_04833_),
    .A2(_04837_),
    .B(_04846_),
    .ZN(_00942_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10181_ (.A1(\u_cpu.cpu.alu.cmp_r ),
    .A2(_02699_),
    .ZN(_04847_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10182_ (.A1(_02699_),
    .A2(_04086_),
    .B(_04847_),
    .ZN(_00943_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10183_ (.I(_02602_),
    .Z(_04848_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10184_ (.I(_04848_),
    .Z(_04849_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10185_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[3] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[2] ),
    .S(_04849_),
    .Z(_04850_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10186_ (.I(_04850_),
    .Z(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10187_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[4] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[3] ),
    .S(_04849_),
    .Z(_04851_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10188_ (.I(_04851_),
    .Z(_00945_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10189_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[5] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[4] ),
    .S(_04849_),
    .Z(_04852_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10190_ (.I(_04852_),
    .Z(_00946_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10191_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[6] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[5] ),
    .S(_04849_),
    .Z(_04853_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10192_ (.I(_04853_),
    .Z(_00947_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10193_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[7] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[6] ),
    .S(_04849_),
    .Z(_04854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10194_ (.I(_04854_),
    .Z(_00948_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10195_ (.I(_04848_),
    .Z(_04855_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10196_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[8] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[7] ),
    .S(_04855_),
    .Z(_04856_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10197_ (.I(_04856_),
    .Z(_00949_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10198_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[9] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[8] ),
    .S(_04855_),
    .Z(_04857_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10199_ (.I(_04857_),
    .Z(_00950_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10200_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[10] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[9] ),
    .S(_04855_),
    .Z(_04858_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10201_ (.I(_04858_),
    .Z(_00951_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10202_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[11] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[10] ),
    .S(_04855_),
    .Z(_04859_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10203_ (.I(_04859_),
    .Z(_00952_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10204_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[12] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[11] ),
    .S(_04855_),
    .Z(_04860_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10205_ (.I(_04860_),
    .Z(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10206_ (.I(_02690_),
    .Z(_04861_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10207_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[13] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[12] ),
    .S(_04861_),
    .Z(_04862_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10208_ (.I(_04862_),
    .Z(_00954_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10209_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[14] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[13] ),
    .S(_04861_),
    .Z(_04863_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10210_ (.I(_04863_),
    .Z(_00955_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10211_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[15] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[14] ),
    .S(_04861_),
    .Z(_04864_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10212_ (.I(_04864_),
    .Z(_00956_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10213_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[16] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[15] ),
    .S(_04861_),
    .Z(_04865_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10214_ (.I(_04865_),
    .Z(_00957_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10215_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[17] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[16] ),
    .S(_04861_),
    .Z(_04866_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10216_ (.I(_04866_),
    .Z(_00958_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10217_ (.I(_02690_),
    .Z(_04867_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10218_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[18] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[17] ),
    .S(_04867_),
    .Z(_04868_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10219_ (.I(_04868_),
    .Z(_00959_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10220_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[19] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[18] ),
    .S(_04867_),
    .Z(_04869_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10221_ (.I(_04869_),
    .Z(_00960_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10222_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[20] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[19] ),
    .S(_04867_),
    .Z(_04870_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10223_ (.I(_04870_),
    .Z(_00961_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10224_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[21] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[20] ),
    .S(_04867_),
    .Z(_04871_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10225_ (.I(_04871_),
    .Z(_00962_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10226_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[22] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[21] ),
    .S(_04867_),
    .Z(_04872_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10227_ (.I(_04872_),
    .Z(_00963_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10228_ (.I(_02690_),
    .Z(_04873_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10229_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[23] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[22] ),
    .S(_04873_),
    .Z(_04874_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10230_ (.I(_04874_),
    .Z(_00964_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10231_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[24] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[23] ),
    .S(_04873_),
    .Z(_04875_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10232_ (.I(_04875_),
    .Z(_00965_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10233_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[25] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[24] ),
    .S(_04873_),
    .Z(_04876_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10234_ (.I(_04876_),
    .Z(_00966_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10235_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[26] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[25] ),
    .S(_04873_),
    .Z(_04877_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10236_ (.I(_04877_),
    .Z(_00967_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10237_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[27] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[26] ),
    .S(_04873_),
    .Z(_04878_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10238_ (.I(_04878_),
    .Z(_00968_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10239_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[28] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[27] ),
    .S(_04848_),
    .Z(_04879_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10240_ (.I(_04879_),
    .Z(_00969_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10241_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[29] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[28] ),
    .S(_04848_),
    .Z(_04880_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10242_ (.I(_04880_),
    .Z(_00970_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10243_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[30] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[29] ),
    .S(_04848_),
    .Z(_04881_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10244_ (.I(_04881_),
    .Z(_00971_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10245_ (.I(\u_arbiter.i_wb_cpu_dbus_adr[31] ),
    .ZN(_04882_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10246_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[30] ),
    .A2(_02691_),
    .ZN(_04883_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10247_ (.A1(_04882_),
    .A2(_02691_),
    .B(_04883_),
    .ZN(_00972_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10248_ (.A1(\u_cpu.cpu.bufreg.i_sh_signed ),
    .A2(_02705_),
    .B(_02691_),
    .ZN(_04884_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10249_ (.A1(_02675_),
    .A2(_02627_),
    .A3(_02686_),
    .B(_02688_),
    .ZN(_04885_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10250_ (.A1(_02689_),
    .A2(_03123_),
    .A3(_04885_),
    .ZN(_04886_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10251_ (.A1(_04882_),
    .A2(_04884_),
    .B1(_04886_),
    .B2(_02691_),
    .ZN(_00973_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10252_ (.A1(\u_cpu.cpu.state.o_cnt_r[0] ),
    .A2(\u_cpu.cpu.state.o_cnt_r[1] ),
    .B(_02565_),
    .C(_03123_),
    .ZN(_04887_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10253_ (.A1(_02690_),
    .A2(_03123_),
    .B(_04887_),
    .ZN(_04888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10254_ (.A1(_01370_),
    .A2(_04888_),
    .ZN(_04889_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10255_ (.A1(_02591_),
    .A2(_04888_),
    .B(_04889_),
    .ZN(_00974_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10256_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[2] ),
    .A2(_02705_),
    .ZN(_04890_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10257_ (.A1(_04886_),
    .A2(_04890_),
    .ZN(_04891_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10258_ (.A1(_04888_),
    .A2(_04891_),
    .ZN(_04892_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10259_ (.A1(_02672_),
    .A2(_04888_),
    .B(_04892_),
    .ZN(_00975_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10260_ (.A1(_03367_),
    .A2(_02921_),
    .ZN(_04893_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10261_ (.I(_04893_),
    .Z(_04894_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10262_ (.I(_04893_),
    .Z(_04895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10263_ (.A1(\u_cpu.rf_ram.memory[30][0] ),
    .A2(_04895_),
    .ZN(_04896_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10264_ (.A1(_04808_),
    .A2(_04894_),
    .B(_04896_),
    .ZN(_00976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10265_ (.A1(\u_cpu.rf_ram.memory[30][1] ),
    .A2(_04895_),
    .ZN(_04897_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10266_ (.A1(_04814_),
    .A2(_04894_),
    .B(_04897_),
    .ZN(_00977_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10267_ (.I(_04893_),
    .Z(_04898_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10268_ (.A1(\u_cpu.rf_ram.memory[30][2] ),
    .A2(_04898_),
    .ZN(_04899_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10269_ (.A1(_04817_),
    .A2(_04894_),
    .B(_04899_),
    .ZN(_00978_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10270_ (.A1(\u_cpu.rf_ram.memory[30][3] ),
    .A2(_04898_),
    .ZN(_04900_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10271_ (.A1(_04821_),
    .A2(_04894_),
    .B(_04900_),
    .ZN(_00979_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10272_ (.A1(\u_cpu.rf_ram.memory[30][4] ),
    .A2(_04898_),
    .ZN(_04901_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10273_ (.A1(_04824_),
    .A2(_04894_),
    .B(_04901_),
    .ZN(_00980_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10274_ (.A1(\u_cpu.rf_ram.memory[30][5] ),
    .A2(_04898_),
    .ZN(_04902_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10275_ (.A1(_04827_),
    .A2(_04895_),
    .B(_04902_),
    .ZN(_00981_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10276_ (.A1(\u_cpu.rf_ram.memory[30][6] ),
    .A2(_04898_),
    .ZN(_04903_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10277_ (.A1(_04830_),
    .A2(_04895_),
    .B(_04903_),
    .ZN(_00982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10278_ (.A1(\u_cpu.rf_ram.memory[30][7] ),
    .A2(_04893_),
    .ZN(_04904_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10279_ (.A1(_04833_),
    .A2(_04895_),
    .B(_04904_),
    .ZN(_00983_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10280_ (.A1(_02528_),
    .A2(_02705_),
    .B(net2),
    .ZN(_04905_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10281_ (.I(_04905_),
    .Z(_04906_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10282_ (.I(_04906_),
    .Z(_04907_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10283_ (.A1(net2),
    .A2(_02696_),
    .ZN(_04908_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10284_ (.I(_04908_),
    .Z(_04909_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10285_ (.I(_04909_),
    .Z(_04910_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10286_ (.A1(_01431_),
    .A2(_04907_),
    .B1(_04910_),
    .B2(\u_arbiter.i_wb_cpu_ibus_adr[1] ),
    .ZN(_04911_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10287_ (.I(_04911_),
    .ZN(_00984_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10288_ (.A1(\u_arbiter.i_wb_cpu_ibus_adr[1] ),
    .A2(_04907_),
    .B1(_04910_),
    .B2(_01444_),
    .ZN(_04912_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10289_ (.I(_04912_),
    .ZN(_00985_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10290_ (.A1(_01444_),
    .A2(_04907_),
    .B1(_04910_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[3] ),
    .ZN(_04913_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10291_ (.I(_04913_),
    .ZN(_00986_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10292_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[3] ),
    .A2(_04907_),
    .B1(_04910_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[4] ),
    .ZN(_04914_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10293_ (.I(_04914_),
    .ZN(_00987_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10294_ (.I(_04906_),
    .Z(_04915_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10295_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[4] ),
    .A2(_04915_),
    .B1(_04910_),
    .B2(_01463_),
    .ZN(_04916_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10296_ (.I(_04916_),
    .ZN(_00988_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10297_ (.I(_04909_),
    .Z(_04917_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10298_ (.A1(_01463_),
    .A2(_04915_),
    .B1(_04917_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[6] ),
    .ZN(_04918_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10299_ (.I(_04918_),
    .ZN(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10300_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[6] ),
    .A2(_04915_),
    .B1(_04917_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[7] ),
    .ZN(_04919_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10301_ (.I(_04919_),
    .ZN(_00990_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10302_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[7] ),
    .A2(_04915_),
    .B1(_04917_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[8] ),
    .ZN(_04920_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10303_ (.I(_04920_),
    .ZN(_00991_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10304_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[8] ),
    .A2(_04915_),
    .B1(_04917_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[9] ),
    .ZN(_04921_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10305_ (.I(_04921_),
    .ZN(_00992_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10306_ (.I(_04905_),
    .Z(_04922_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10307_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[9] ),
    .A2(_04922_),
    .B1(_04917_),
    .B2(_01484_),
    .ZN(_04923_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10308_ (.I(_04923_),
    .ZN(_00993_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10309_ (.I(_04909_),
    .Z(_04924_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10310_ (.A1(_01484_),
    .A2(_04922_),
    .B1(_04924_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[11] ),
    .ZN(_04925_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10311_ (.I(_04925_),
    .ZN(_00994_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10312_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[11] ),
    .A2(_04922_),
    .B1(_04924_),
    .B2(_01495_),
    .ZN(_04926_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10313_ (.I(_04926_),
    .ZN(_00995_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10314_ (.A1(_01495_),
    .A2(_04922_),
    .B1(_04924_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[13] ),
    .ZN(_04927_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10315_ (.I(_04927_),
    .ZN(_00996_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10316_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[13] ),
    .A2(_04922_),
    .B1(_04924_),
    .B2(_01502_),
    .ZN(_04928_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10317_ (.I(_04928_),
    .ZN(_00997_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10318_ (.I(_04905_),
    .Z(_04929_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10319_ (.A1(_01502_),
    .A2(_04929_),
    .B1(_04924_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[15] ),
    .ZN(_04930_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10320_ (.I(_04930_),
    .ZN(_00998_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10321_ (.I(_04908_),
    .Z(_04931_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10322_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[15] ),
    .A2(_04929_),
    .B1(_04931_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[16] ),
    .ZN(_04932_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10323_ (.I(_04932_),
    .ZN(_00999_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10324_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[16] ),
    .A2(_04929_),
    .B1(_04931_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[17] ),
    .ZN(_04933_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10325_ (.I(_04933_),
    .ZN(_01000_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10326_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[17] ),
    .A2(_04929_),
    .B1(_04931_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[18] ),
    .ZN(_04934_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10327_ (.I(_04934_),
    .ZN(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10328_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[18] ),
    .A2(_04929_),
    .B1(_04931_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[19] ),
    .ZN(_04935_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10329_ (.I(_04935_),
    .ZN(_01002_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10330_ (.I(_04905_),
    .Z(_04936_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10331_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[19] ),
    .A2(_04936_),
    .B1(_04931_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[20] ),
    .ZN(_04937_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10332_ (.I(_04937_),
    .ZN(_01003_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10333_ (.I(_04908_),
    .Z(_04938_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10334_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[20] ),
    .A2(_04936_),
    .B1(_04938_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[21] ),
    .ZN(_04939_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10335_ (.I(_04939_),
    .ZN(_01004_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10336_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[21] ),
    .A2(_04936_),
    .B1(_04938_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[22] ),
    .ZN(_04940_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10337_ (.I(_04940_),
    .ZN(_01005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10338_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[22] ),
    .A2(_04936_),
    .B1(_04938_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[23] ),
    .ZN(_04941_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10339_ (.I(_04941_),
    .ZN(_01006_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10340_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[23] ),
    .A2(_04936_),
    .B1(_04938_),
    .B2(_01537_),
    .ZN(_04942_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10341_ (.I(_04942_),
    .ZN(_01007_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10342_ (.I(_04905_),
    .Z(_04943_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10343_ (.A1(_01537_),
    .A2(_04943_),
    .B1(_04938_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[25] ),
    .ZN(_04944_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10344_ (.I(_04944_),
    .ZN(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10345_ (.I(_04908_),
    .Z(_04945_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10346_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[25] ),
    .A2(_04943_),
    .B1(_04945_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[26] ),
    .ZN(_04946_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10347_ (.I(_04946_),
    .ZN(_01009_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10348_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[26] ),
    .A2(_04943_),
    .B1(_04945_),
    .B2(_01547_),
    .ZN(_04947_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10349_ (.I(_04947_),
    .ZN(_01010_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10350_ (.A1(_01547_),
    .A2(_04943_),
    .B1(_04945_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[28] ),
    .ZN(_04948_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10351_ (.I(_04948_),
    .ZN(_01011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10352_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[28] ),
    .A2(_04943_),
    .B1(_04945_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[29] ),
    .ZN(_04949_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10353_ (.I(_04949_),
    .ZN(_01012_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10354_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[29] ),
    .A2(_04906_),
    .B1(_04945_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[30] ),
    .ZN(_04950_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10355_ (.I(_04950_),
    .ZN(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10356_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[30] ),
    .A2(_04906_),
    .B1(_04909_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[31] ),
    .ZN(_04951_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10357_ (.I(_04951_),
    .ZN(_01014_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10358_ (.A1(_02571_),
    .A2(_01412_),
    .A3(_01379_),
    .ZN(_04952_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10359_ (.A1(_04952_),
    .A2(_02579_),
    .ZN(_04953_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10360_ (.I0(_02612_),
    .I1(_02640_),
    .S(\u_cpu.cpu.ctrl.i_jump ),
    .Z(_04954_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10361_ (.A1(_02545_),
    .A2(_02586_),
    .B(_04953_),
    .ZN(_04955_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10362_ (.A1(_04953_),
    .A2(_04954_),
    .B(_04955_),
    .ZN(_04956_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10363_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[31] ),
    .A2(_04906_),
    .B1(_04909_),
    .B2(_04956_),
    .ZN(_04957_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10364_ (.I(_04957_),
    .ZN(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10365_ (.A1(_02700_),
    .A2(_02729_),
    .A3(_02847_),
    .ZN(_04958_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10366_ (.I(_04958_),
    .Z(_04959_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10367_ (.A1(_02966_),
    .A2(_04959_),
    .ZN(_04960_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10368_ (.I(_04960_),
    .Z(_04961_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10369_ (.I(_04960_),
    .Z(_04962_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10370_ (.A1(\u_cpu.rf_ram.memory[109][0] ),
    .A2(_04962_),
    .ZN(_04963_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10371_ (.A1(_04808_),
    .A2(_04961_),
    .B(_04963_),
    .ZN(_01016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10372_ (.A1(\u_cpu.rf_ram.memory[109][1] ),
    .A2(_04962_),
    .ZN(_04964_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10373_ (.A1(_04814_),
    .A2(_04961_),
    .B(_04964_),
    .ZN(_01017_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10374_ (.I(_04960_),
    .Z(_04965_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10375_ (.A1(\u_cpu.rf_ram.memory[109][2] ),
    .A2(_04965_),
    .ZN(_04966_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10376_ (.A1(_04817_),
    .A2(_04961_),
    .B(_04966_),
    .ZN(_01018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10377_ (.A1(\u_cpu.rf_ram.memory[109][3] ),
    .A2(_04965_),
    .ZN(_04967_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10378_ (.A1(_04821_),
    .A2(_04961_),
    .B(_04967_),
    .ZN(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10379_ (.A1(\u_cpu.rf_ram.memory[109][4] ),
    .A2(_04965_),
    .ZN(_04968_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10380_ (.A1(_04824_),
    .A2(_04961_),
    .B(_04968_),
    .ZN(_01020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10381_ (.A1(\u_cpu.rf_ram.memory[109][5] ),
    .A2(_04965_),
    .ZN(_04969_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10382_ (.A1(_04827_),
    .A2(_04962_),
    .B(_04969_),
    .ZN(_01021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10383_ (.A1(\u_cpu.rf_ram.memory[109][6] ),
    .A2(_04965_),
    .ZN(_04970_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10384_ (.A1(_04830_),
    .A2(_04962_),
    .B(_04970_),
    .ZN(_01022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10385_ (.A1(\u_cpu.rf_ram.memory[109][7] ),
    .A2(_04960_),
    .ZN(_04971_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10386_ (.A1(_04833_),
    .A2(_04962_),
    .B(_04971_),
    .ZN(_01023_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10387_ (.A1(_03870_),
    .A2(_03310_),
    .ZN(_04972_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10388_ (.I(_04972_),
    .Z(_04973_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10389_ (.I0(_04184_),
    .I1(\u_cpu.rf_ram.memory[3][0] ),
    .S(_04973_),
    .Z(_04974_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10390_ (.I(_04974_),
    .Z(_01024_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10391_ (.I0(_04188_),
    .I1(\u_cpu.rf_ram.memory[3][1] ),
    .S(_04973_),
    .Z(_04975_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10392_ (.I(_04975_),
    .Z(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10393_ (.I0(_04190_),
    .I1(\u_cpu.rf_ram.memory[3][2] ),
    .S(_04973_),
    .Z(_04976_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10394_ (.I(_04976_),
    .Z(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10395_ (.I0(_04192_),
    .I1(\u_cpu.rf_ram.memory[3][3] ),
    .S(_04973_),
    .Z(_04977_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10396_ (.I(_04977_),
    .Z(_01027_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10397_ (.I0(_04194_),
    .I1(\u_cpu.rf_ram.memory[3][4] ),
    .S(_04973_),
    .Z(_04978_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10398_ (.I(_04978_),
    .Z(_01028_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10399_ (.I0(_04196_),
    .I1(\u_cpu.rf_ram.memory[3][5] ),
    .S(_04972_),
    .Z(_04979_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10400_ (.I(_04979_),
    .Z(_01029_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10401_ (.I0(_04198_),
    .I1(\u_cpu.rf_ram.memory[3][6] ),
    .S(_04972_),
    .Z(_04980_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10402_ (.I(_04980_),
    .Z(_01030_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10403_ (.I0(_04200_),
    .I1(\u_cpu.rf_ram.memory[3][7] ),
    .S(_04972_),
    .Z(_04981_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10404_ (.I(_04981_),
    .Z(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10405_ (.A1(_02723_),
    .A2(_02850_),
    .ZN(_04982_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10406_ (.I(_04982_),
    .Z(_04983_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10407_ (.I0(_04184_),
    .I1(\u_cpu.rf_ram.memory[2][0] ),
    .S(_04983_),
    .Z(_04984_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10408_ (.I(_04984_),
    .Z(_01032_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10409_ (.I0(_04188_),
    .I1(\u_cpu.rf_ram.memory[2][1] ),
    .S(_04983_),
    .Z(_04985_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10410_ (.I(_04985_),
    .Z(_01033_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10411_ (.I0(_04190_),
    .I1(\u_cpu.rf_ram.memory[2][2] ),
    .S(_04983_),
    .Z(_04986_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10412_ (.I(_04986_),
    .Z(_01034_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10413_ (.I0(_04192_),
    .I1(\u_cpu.rf_ram.memory[2][3] ),
    .S(_04983_),
    .Z(_04987_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10414_ (.I(_04987_),
    .Z(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10415_ (.I0(_04194_),
    .I1(\u_cpu.rf_ram.memory[2][4] ),
    .S(_04983_),
    .Z(_04988_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10416_ (.I(_04988_),
    .Z(_01036_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10417_ (.I0(_04196_),
    .I1(\u_cpu.rf_ram.memory[2][5] ),
    .S(_04982_),
    .Z(_04989_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10418_ (.I(_04989_),
    .Z(_01037_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10419_ (.I0(_04198_),
    .I1(\u_cpu.rf_ram.memory[2][6] ),
    .S(_04982_),
    .Z(_04990_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10420_ (.I(_04990_),
    .Z(_01038_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10421_ (.I0(_04200_),
    .I1(\u_cpu.rf_ram.memory[2][7] ),
    .S(_04982_),
    .Z(_04991_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10422_ (.I(_04991_),
    .Z(_01039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10423_ (.A1(_04091_),
    .A2(_02967_),
    .ZN(_04992_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10424_ (.I(_04992_),
    .Z(_04993_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10425_ (.I(_04992_),
    .Z(_04994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10426_ (.A1(\u_cpu.rf_ram.memory[93][0] ),
    .A2(_04994_),
    .ZN(_04995_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10427_ (.A1(_04808_),
    .A2(_04993_),
    .B(_04995_),
    .ZN(_01040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10428_ (.A1(\u_cpu.rf_ram.memory[93][1] ),
    .A2(_04994_),
    .ZN(_04996_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10429_ (.A1(_04814_),
    .A2(_04993_),
    .B(_04996_),
    .ZN(_01041_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10430_ (.I(_04992_),
    .Z(_04997_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10431_ (.A1(\u_cpu.rf_ram.memory[93][2] ),
    .A2(_04997_),
    .ZN(_04998_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10432_ (.A1(_04817_),
    .A2(_04993_),
    .B(_04998_),
    .ZN(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10433_ (.A1(\u_cpu.rf_ram.memory[93][3] ),
    .A2(_04997_),
    .ZN(_04999_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10434_ (.A1(_04821_),
    .A2(_04993_),
    .B(_04999_),
    .ZN(_01043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10435_ (.A1(\u_cpu.rf_ram.memory[93][4] ),
    .A2(_04997_),
    .ZN(_05000_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10436_ (.A1(_04824_),
    .A2(_04993_),
    .B(_05000_),
    .ZN(_01044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10437_ (.A1(\u_cpu.rf_ram.memory[93][5] ),
    .A2(_04997_),
    .ZN(_05001_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10438_ (.A1(_04827_),
    .A2(_04994_),
    .B(_05001_),
    .ZN(_01045_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10439_ (.A1(\u_cpu.rf_ram.memory[93][6] ),
    .A2(_04997_),
    .ZN(_05002_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10440_ (.A1(_04830_),
    .A2(_04994_),
    .B(_05002_),
    .ZN(_01046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10441_ (.A1(\u_cpu.rf_ram.memory[93][7] ),
    .A2(_04992_),
    .ZN(_05003_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10442_ (.A1(_04833_),
    .A2(_04994_),
    .B(_05003_),
    .ZN(_01047_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10443_ (.A1(_02674_),
    .A2(_02704_),
    .ZN(_05004_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10444_ (.A1(_03118_),
    .A2(_05004_),
    .ZN(_05005_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10445_ (.I(_05005_),
    .Z(_05006_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10446_ (.A1(\u_cpu.cpu.immdec.imm11_7[1] ),
    .A2(_04636_),
    .B(_05005_),
    .ZN(_05007_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10447_ (.A1(_02535_),
    .A2(_05006_),
    .B1(_05007_),
    .B2(_04732_),
    .ZN(_01048_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10448_ (.A1(_04566_),
    .A2(_04503_),
    .B(_04602_),
    .ZN(_05008_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10449_ (.A1(_04562_),
    .A2(_04700_),
    .A3(_05008_),
    .ZN(_05009_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10450_ (.A1(_04763_),
    .A2(_05009_),
    .B(_04560_),
    .ZN(_05010_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _10451_ (.A1(_04407_),
    .A2(_04518_),
    .A3(_04722_),
    .B1(_05010_),
    .B2(_04469_),
    .ZN(_05011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10452_ (.A1(_04468_),
    .A2(_04510_),
    .B1(_04652_),
    .B2(_04680_),
    .ZN(_05012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10453_ (.A1(_04560_),
    .A2(_05012_),
    .ZN(_05013_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10454_ (.A1(_04398_),
    .A2(_05011_),
    .A3(_05013_),
    .ZN(_05014_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10455_ (.I0(\u_cpu.cpu.immdec.imm11_7[1] ),
    .I1(_02700_),
    .S(_05004_),
    .Z(_05015_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10456_ (.A1(_04680_),
    .A2(_04500_),
    .B1(_05015_),
    .B2(_04482_),
    .ZN(_05016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10457_ (.A1(_05014_),
    .A2(_05016_),
    .ZN(_01049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10458_ (.A1(_04497_),
    .A2(_04509_),
    .ZN(_05017_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _10459_ (.A1(_04692_),
    .A2(_04433_),
    .B1(_04491_),
    .B2(_04514_),
    .C(_05017_),
    .ZN(_05018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10460_ (.A1(_04401_),
    .A2(_04520_),
    .ZN(_05019_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10461_ (.A1(_04492_),
    .A2(_05019_),
    .B(_04700_),
    .C(_04581_),
    .ZN(_05020_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10462_ (.A1(_04444_),
    .A2(_05018_),
    .B1(_05020_),
    .B2(_04747_),
    .ZN(_05021_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10463_ (.A1(_04494_),
    .A2(_05021_),
    .ZN(_05022_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10464_ (.A1(_02701_),
    .A2(_04630_),
    .B(_05022_),
    .ZN(_05023_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10465_ (.A1(_04518_),
    .A2(_04434_),
    .ZN(_05024_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10466_ (.A1(_04446_),
    .A2(_05024_),
    .ZN(_05025_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10467_ (.A1(_04692_),
    .A2(_05025_),
    .ZN(_05026_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10468_ (.A1(_02700_),
    .A2(_05006_),
    .B1(_05026_),
    .B2(_04516_),
    .ZN(_05027_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10469_ (.A1(_05006_),
    .A2(_05023_),
    .B(_05027_),
    .ZN(_01050_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10470_ (.A1(_04419_),
    .A2(_04452_),
    .B(_05025_),
    .C(_04582_),
    .ZN(_05028_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10471_ (.A1(_04510_),
    .A2(_04560_),
    .B1(_05028_),
    .B2(_04701_),
    .ZN(_05029_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10472_ (.A1(_04525_),
    .A2(_04613_),
    .B(_05029_),
    .ZN(_05030_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10473_ (.A1(_02701_),
    .A2(_05004_),
    .ZN(_05031_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10474_ (.A1(_02787_),
    .A2(_05004_),
    .B(_05031_),
    .ZN(_05032_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10475_ (.I0(_05030_),
    .I1(_05032_),
    .S(_04466_),
    .Z(_05033_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10476_ (.I(_05033_),
    .Z(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10477_ (.A1(_04545_),
    .A2(_04453_),
    .ZN(_05034_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10478_ (.A1(_04567_),
    .A2(_05034_),
    .B(_04487_),
    .C(_04575_),
    .ZN(_05035_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10479_ (.A1(_04493_),
    .A2(_04491_),
    .A3(_05035_),
    .ZN(_05036_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10480_ (.A1(_04516_),
    .A2(_04650_),
    .A3(_05036_),
    .ZN(_05037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10481_ (.A1(\u_cpu.cpu.immdec.imm30_25[0] ),
    .A2(_04630_),
    .B(_05006_),
    .ZN(_05038_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10482_ (.A1(_02787_),
    .A2(_05006_),
    .B1(_05037_),
    .B2(_05038_),
    .ZN(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10483_ (.I(_04807_),
    .Z(_05039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10484_ (.A1(_02803_),
    .A2(_04959_),
    .ZN(_05040_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10485_ (.I(_05040_),
    .Z(_05041_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10486_ (.I(_05040_),
    .Z(_05042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10487_ (.A1(\u_cpu.rf_ram.memory[97][0] ),
    .A2(_05042_),
    .ZN(_05043_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10488_ (.A1(_05039_),
    .A2(_05041_),
    .B(_05043_),
    .ZN(_01053_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10489_ (.I(_04813_),
    .Z(_05044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10490_ (.A1(\u_cpu.rf_ram.memory[97][1] ),
    .A2(_05042_),
    .ZN(_05045_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10491_ (.A1(_05044_),
    .A2(_05041_),
    .B(_05045_),
    .ZN(_01054_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10492_ (.I(_04816_),
    .Z(_05046_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10493_ (.I(_05040_),
    .Z(_05047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10494_ (.A1(\u_cpu.rf_ram.memory[97][2] ),
    .A2(_05047_),
    .ZN(_05048_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10495_ (.A1(_05046_),
    .A2(_05041_),
    .B(_05048_),
    .ZN(_01055_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10496_ (.I(_04820_),
    .Z(_05049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10497_ (.A1(\u_cpu.rf_ram.memory[97][3] ),
    .A2(_05047_),
    .ZN(_05050_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10498_ (.A1(_05049_),
    .A2(_05041_),
    .B(_05050_),
    .ZN(_01056_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10499_ (.I(_04823_),
    .Z(_05051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10500_ (.A1(\u_cpu.rf_ram.memory[97][4] ),
    .A2(_05047_),
    .ZN(_05052_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10501_ (.A1(_05051_),
    .A2(_05041_),
    .B(_05052_),
    .ZN(_01057_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10502_ (.I(_04826_),
    .Z(_05053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10503_ (.A1(\u_cpu.rf_ram.memory[97][5] ),
    .A2(_05047_),
    .ZN(_05054_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10504_ (.A1(_05053_),
    .A2(_05042_),
    .B(_05054_),
    .ZN(_01058_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10505_ (.I(_04829_),
    .Z(_05055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10506_ (.A1(\u_cpu.rf_ram.memory[97][6] ),
    .A2(_05047_),
    .ZN(_05056_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10507_ (.A1(_05055_),
    .A2(_05042_),
    .B(_05056_),
    .ZN(_01059_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10508_ (.I(_04832_),
    .Z(_05057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10509_ (.A1(\u_cpu.rf_ram.memory[97][7] ),
    .A2(_05040_),
    .ZN(_05058_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10510_ (.A1(_05057_),
    .A2(_05042_),
    .B(_05058_),
    .ZN(_01060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10511_ (.A1(_04091_),
    .A2(_02921_),
    .ZN(_05059_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10512_ (.I(_05059_),
    .Z(_05060_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10513_ (.I(_05059_),
    .Z(_05061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10514_ (.A1(\u_cpu.rf_ram.memory[94][0] ),
    .A2(_05061_),
    .ZN(_05062_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10515_ (.A1(_05039_),
    .A2(_05060_),
    .B(_05062_),
    .ZN(_01061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10516_ (.A1(\u_cpu.rf_ram.memory[94][1] ),
    .A2(_05061_),
    .ZN(_05063_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10517_ (.A1(_05044_),
    .A2(_05060_),
    .B(_05063_),
    .ZN(_01062_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10518_ (.I(_05059_),
    .Z(_05064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10519_ (.A1(\u_cpu.rf_ram.memory[94][2] ),
    .A2(_05064_),
    .ZN(_05065_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10520_ (.A1(_05046_),
    .A2(_05060_),
    .B(_05065_),
    .ZN(_01063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10521_ (.A1(\u_cpu.rf_ram.memory[94][3] ),
    .A2(_05064_),
    .ZN(_05066_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10522_ (.A1(_05049_),
    .A2(_05060_),
    .B(_05066_),
    .ZN(_01064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10523_ (.A1(\u_cpu.rf_ram.memory[94][4] ),
    .A2(_05064_),
    .ZN(_05067_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10524_ (.A1(_05051_),
    .A2(_05060_),
    .B(_05067_),
    .ZN(_01065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10525_ (.A1(\u_cpu.rf_ram.memory[94][5] ),
    .A2(_05064_),
    .ZN(_05068_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10526_ (.A1(_05053_),
    .A2(_05061_),
    .B(_05068_),
    .ZN(_01066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10527_ (.A1(\u_cpu.rf_ram.memory[94][6] ),
    .A2(_05064_),
    .ZN(_05069_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10528_ (.A1(_05055_),
    .A2(_05061_),
    .B(_05069_),
    .ZN(_01067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10529_ (.A1(\u_cpu.rf_ram.memory[94][7] ),
    .A2(_05059_),
    .ZN(_05070_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10530_ (.A1(_05057_),
    .A2(_05061_),
    .B(_05070_),
    .ZN(_01068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10531_ (.A1(_04091_),
    .A2(_03062_),
    .ZN(_05071_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10532_ (.I(_05071_),
    .Z(_05072_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10533_ (.I(_05071_),
    .Z(_05073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10534_ (.A1(\u_cpu.rf_ram.memory[95][0] ),
    .A2(_05073_),
    .ZN(_05074_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10535_ (.A1(_05039_),
    .A2(_05072_),
    .B(_05074_),
    .ZN(_01069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10536_ (.A1(\u_cpu.rf_ram.memory[95][1] ),
    .A2(_05073_),
    .ZN(_05075_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10537_ (.A1(_05044_),
    .A2(_05072_),
    .B(_05075_),
    .ZN(_01070_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10538_ (.I(_05071_),
    .Z(_05076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10539_ (.A1(\u_cpu.rf_ram.memory[95][2] ),
    .A2(_05076_),
    .ZN(_05077_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10540_ (.A1(_05046_),
    .A2(_05072_),
    .B(_05077_),
    .ZN(_01071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10541_ (.A1(\u_cpu.rf_ram.memory[95][3] ),
    .A2(_05076_),
    .ZN(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10542_ (.A1(_05049_),
    .A2(_05072_),
    .B(_05078_),
    .ZN(_01072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10543_ (.A1(\u_cpu.rf_ram.memory[95][4] ),
    .A2(_05076_),
    .ZN(_05079_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10544_ (.A1(_05051_),
    .A2(_05072_),
    .B(_05079_),
    .ZN(_01073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10545_ (.A1(\u_cpu.rf_ram.memory[95][5] ),
    .A2(_05076_),
    .ZN(_05080_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10546_ (.A1(_05053_),
    .A2(_05073_),
    .B(_05080_),
    .ZN(_01074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10547_ (.A1(\u_cpu.rf_ram.memory[95][6] ),
    .A2(_05076_),
    .ZN(_05081_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10548_ (.A1(_05055_),
    .A2(_05073_),
    .B(_05081_),
    .ZN(_01075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10549_ (.A1(\u_cpu.rf_ram.memory[95][7] ),
    .A2(_05071_),
    .ZN(_05082_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10550_ (.A1(_05057_),
    .A2(_05073_),
    .B(_05082_),
    .ZN(_01076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10551_ (.A1(_02890_),
    .A2(_04959_),
    .ZN(_05083_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10552_ (.I(_05083_),
    .Z(_05084_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10553_ (.I(_05083_),
    .Z(_05085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10554_ (.A1(\u_cpu.rf_ram.memory[96][0] ),
    .A2(_05085_),
    .ZN(_05086_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10555_ (.A1(_05039_),
    .A2(_05084_),
    .B(_05086_),
    .ZN(_01077_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10556_ (.A1(\u_cpu.rf_ram.memory[96][1] ),
    .A2(_05085_),
    .ZN(_05087_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10557_ (.A1(_05044_),
    .A2(_05084_),
    .B(_05087_),
    .ZN(_01078_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10558_ (.I(_05083_),
    .Z(_05088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10559_ (.A1(\u_cpu.rf_ram.memory[96][2] ),
    .A2(_05088_),
    .ZN(_05089_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10560_ (.A1(_05046_),
    .A2(_05084_),
    .B(_05089_),
    .ZN(_01079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10561_ (.A1(\u_cpu.rf_ram.memory[96][3] ),
    .A2(_05088_),
    .ZN(_05090_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10562_ (.A1(_05049_),
    .A2(_05084_),
    .B(_05090_),
    .ZN(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10563_ (.A1(\u_cpu.rf_ram.memory[96][4] ),
    .A2(_05088_),
    .ZN(_05091_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10564_ (.A1(_05051_),
    .A2(_05084_),
    .B(_05091_),
    .ZN(_01081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10565_ (.A1(\u_cpu.rf_ram.memory[96][5] ),
    .A2(_05088_),
    .ZN(_05092_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10566_ (.A1(_05053_),
    .A2(_05085_),
    .B(_05092_),
    .ZN(_01082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10567_ (.A1(\u_cpu.rf_ram.memory[96][6] ),
    .A2(_05088_),
    .ZN(_05093_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10568_ (.A1(_05055_),
    .A2(_05085_),
    .B(_05093_),
    .ZN(_01083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10569_ (.A1(\u_cpu.rf_ram.memory[96][7] ),
    .A2(_05083_),
    .ZN(_05094_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10570_ (.A1(_05057_),
    .A2(_05085_),
    .B(_05094_),
    .ZN(_01084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10571_ (.A1(\u_cpu.cpu.bufreg.i_sh_signed ),
    .A2(_04467_),
    .ZN(_05095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10572_ (.A1(_04713_),
    .A2(_05095_),
    .ZN(_01085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10573_ (.A1(\u_arbiter.i_wb_cpu_ack ),
    .A2(\u_arbiter.o_wb_cpu_adr[1] ),
    .ZN(_05096_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10574_ (.A1(_01443_),
    .A2(_05096_),
    .Z(_05097_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10575_ (.A1(_03112_),
    .A2(_05097_),
    .ZN(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10576_ (.I(_02789_),
    .Z(_05098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10577_ (.A1(_05098_),
    .A2(_02982_),
    .ZN(_05099_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10578_ (.I(_05099_),
    .Z(_05100_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10579_ (.I(_05099_),
    .Z(_05101_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10580_ (.A1(\u_cpu.rf_ram.memory[28][0] ),
    .A2(_05101_),
    .ZN(_05102_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10581_ (.A1(_05039_),
    .A2(_05100_),
    .B(_05102_),
    .ZN(_01087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10582_ (.A1(\u_cpu.rf_ram.memory[28][1] ),
    .A2(_05101_),
    .ZN(_05103_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10583_ (.A1(_05044_),
    .A2(_05100_),
    .B(_05103_),
    .ZN(_01088_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10584_ (.I(_05099_),
    .Z(_05104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10585_ (.A1(\u_cpu.rf_ram.memory[28][2] ),
    .A2(_05104_),
    .ZN(_05105_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10586_ (.A1(_05046_),
    .A2(_05100_),
    .B(_05105_),
    .ZN(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10587_ (.A1(\u_cpu.rf_ram.memory[28][3] ),
    .A2(_05104_),
    .ZN(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10588_ (.A1(_05049_),
    .A2(_05100_),
    .B(_05106_),
    .ZN(_01090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10589_ (.A1(\u_cpu.rf_ram.memory[28][4] ),
    .A2(_05104_),
    .ZN(_05107_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10590_ (.A1(_05051_),
    .A2(_05100_),
    .B(_05107_),
    .ZN(_01091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10591_ (.A1(\u_cpu.rf_ram.memory[28][5] ),
    .A2(_05104_),
    .ZN(_05108_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10592_ (.A1(_05053_),
    .A2(_05101_),
    .B(_05108_),
    .ZN(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10593_ (.A1(\u_cpu.rf_ram.memory[28][6] ),
    .A2(_05104_),
    .ZN(_05109_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10594_ (.A1(_05055_),
    .A2(_05101_),
    .B(_05109_),
    .ZN(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10595_ (.A1(\u_cpu.rf_ram.memory[28][7] ),
    .A2(_05099_),
    .ZN(_05110_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10596_ (.A1(_05057_),
    .A2(_05101_),
    .B(_05110_),
    .ZN(_01094_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10597_ (.I(_03116_),
    .Z(_05111_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10598_ (.I0(\u_arbiter.i_wb_cpu_rdt[16] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ),
    .S(_05111_),
    .Z(_05112_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10599_ (.I(_05112_),
    .Z(_01095_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10600_ (.I0(\u_arbiter.i_wb_cpu_rdt[17] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ),
    .S(_05111_),
    .Z(_05113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10601_ (.I(_05113_),
    .Z(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10602_ (.I0(\u_arbiter.i_wb_cpu_rdt[18] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[2] ),
    .S(_05111_),
    .Z(_05114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10603_ (.I(_05114_),
    .Z(_01097_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10604_ (.I0(\u_arbiter.i_wb_cpu_rdt[19] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[3] ),
    .S(_05111_),
    .Z(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10605_ (.I(_05115_),
    .Z(_01098_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10606_ (.I0(\u_arbiter.i_wb_cpu_rdt[20] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ),
    .S(_05111_),
    .Z(_05116_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10607_ (.I(_05116_),
    .Z(_01099_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10608_ (.I(_03116_),
    .Z(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10609_ (.I0(\u_arbiter.i_wb_cpu_rdt[21] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ),
    .S(_05117_),
    .Z(_05118_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10610_ (.I(_05118_),
    .Z(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10611_ (.I0(\u_arbiter.i_wb_cpu_rdt[22] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ),
    .S(_05117_),
    .Z(_05119_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10612_ (.I(_05119_),
    .Z(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10613_ (.I0(\u_arbiter.i_wb_cpu_rdt[23] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ),
    .S(_05117_),
    .Z(_05120_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10614_ (.I(_05120_),
    .Z(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10615_ (.I0(\u_arbiter.i_wb_cpu_rdt[24] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ),
    .S(_05117_),
    .Z(_05121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10616_ (.I(_05121_),
    .Z(_01103_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10617_ (.I0(\u_arbiter.i_wb_cpu_rdt[25] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ),
    .S(_05117_),
    .Z(_05122_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10618_ (.I(_05122_),
    .Z(_01104_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10619_ (.I(_03116_),
    .Z(_05123_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10620_ (.I0(\u_arbiter.i_wb_cpu_rdt[26] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[10] ),
    .S(_05123_),
    .Z(_05124_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10621_ (.I(_05124_),
    .Z(_01105_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10622_ (.I0(\u_arbiter.i_wb_cpu_rdt[27] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[11] ),
    .S(_05123_),
    .Z(_05125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10623_ (.I(_05125_),
    .Z(_01106_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10624_ (.I0(\u_arbiter.i_wb_cpu_rdt[28] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ),
    .S(_05123_),
    .Z(_05126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10625_ (.I(_05126_),
    .Z(_01107_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10626_ (.I0(\u_arbiter.i_wb_cpu_rdt[29] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ),
    .S(_05123_),
    .Z(_05127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10627_ (.I(_05127_),
    .Z(_01108_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10628_ (.I0(\u_arbiter.i_wb_cpu_rdt[30] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ),
    .S(_05123_),
    .Z(_05128_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10629_ (.I(_05128_),
    .Z(_01109_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10630_ (.I0(\u_arbiter.i_wb_cpu_rdt[31] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ),
    .S(_03116_),
    .Z(_05129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10631_ (.I(_05129_),
    .Z(_01110_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10632_ (.I(_04807_),
    .Z(_05130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10633_ (.A1(_02785_),
    .A2(_04959_),
    .ZN(_05131_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10634_ (.I(_05131_),
    .Z(_05132_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10635_ (.I(_05131_),
    .Z(_05133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10636_ (.A1(\u_cpu.rf_ram.memory[101][0] ),
    .A2(_05133_),
    .ZN(_05134_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10637_ (.A1(_05130_),
    .A2(_05132_),
    .B(_05134_),
    .ZN(_01111_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10638_ (.I(_04813_),
    .Z(_05135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10639_ (.A1(\u_cpu.rf_ram.memory[101][1] ),
    .A2(_05133_),
    .ZN(_05136_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10640_ (.A1(_05135_),
    .A2(_05132_),
    .B(_05136_),
    .ZN(_01112_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10641_ (.I(_04816_),
    .Z(_05137_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10642_ (.I(_05131_),
    .Z(_05138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10643_ (.A1(\u_cpu.rf_ram.memory[101][2] ),
    .A2(_05138_),
    .ZN(_05139_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10644_ (.A1(_05137_),
    .A2(_05132_),
    .B(_05139_),
    .ZN(_01113_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10645_ (.I(_04820_),
    .Z(_05140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10646_ (.A1(\u_cpu.rf_ram.memory[101][3] ),
    .A2(_05138_),
    .ZN(_05141_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10647_ (.A1(_05140_),
    .A2(_05132_),
    .B(_05141_),
    .ZN(_01114_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10648_ (.I(_04823_),
    .Z(_05142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10649_ (.A1(\u_cpu.rf_ram.memory[101][4] ),
    .A2(_05138_),
    .ZN(_05143_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10650_ (.A1(_05142_),
    .A2(_05132_),
    .B(_05143_),
    .ZN(_01115_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10651_ (.I(_04826_),
    .Z(_05144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10652_ (.A1(\u_cpu.rf_ram.memory[101][5] ),
    .A2(_05138_),
    .ZN(_05145_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10653_ (.A1(_05144_),
    .A2(_05133_),
    .B(_05145_),
    .ZN(_01116_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10654_ (.I(_04829_),
    .Z(_05146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10655_ (.A1(\u_cpu.rf_ram.memory[101][6] ),
    .A2(_05138_),
    .ZN(_05147_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10656_ (.A1(_05146_),
    .A2(_05133_),
    .B(_05147_),
    .ZN(_01117_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10657_ (.I(_04832_),
    .Z(_05148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10658_ (.A1(\u_cpu.rf_ram.memory[101][7] ),
    .A2(_05131_),
    .ZN(_05149_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10659_ (.A1(_05148_),
    .A2(_05133_),
    .B(_05149_),
    .ZN(_01118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10660_ (.A1(_03286_),
    .A2(_04959_),
    .ZN(_05150_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10661_ (.I(_05150_),
    .Z(_05151_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10662_ (.I(_05150_),
    .Z(_05152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10663_ (.A1(\u_cpu.rf_ram.memory[102][0] ),
    .A2(_05152_),
    .ZN(_05153_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10664_ (.A1(_05130_),
    .A2(_05151_),
    .B(_05153_),
    .ZN(_01119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10665_ (.A1(\u_cpu.rf_ram.memory[102][1] ),
    .A2(_05152_),
    .ZN(_05154_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10666_ (.A1(_05135_),
    .A2(_05151_),
    .B(_05154_),
    .ZN(_01120_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10667_ (.I(_05150_),
    .Z(_05155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10668_ (.A1(\u_cpu.rf_ram.memory[102][2] ),
    .A2(_05155_),
    .ZN(_05156_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10669_ (.A1(_05137_),
    .A2(_05151_),
    .B(_05156_),
    .ZN(_01121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10670_ (.A1(\u_cpu.rf_ram.memory[102][3] ),
    .A2(_05155_),
    .ZN(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10671_ (.A1(_05140_),
    .A2(_05151_),
    .B(_05157_),
    .ZN(_01122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10672_ (.A1(\u_cpu.rf_ram.memory[102][4] ),
    .A2(_05155_),
    .ZN(_05158_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10673_ (.A1(_05142_),
    .A2(_05151_),
    .B(_05158_),
    .ZN(_01123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10674_ (.A1(\u_cpu.rf_ram.memory[102][5] ),
    .A2(_05155_),
    .ZN(_05159_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10675_ (.A1(_05144_),
    .A2(_05152_),
    .B(_05159_),
    .ZN(_01124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10676_ (.A1(\u_cpu.rf_ram.memory[102][6] ),
    .A2(_05155_),
    .ZN(_05160_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10677_ (.A1(_05146_),
    .A2(_05152_),
    .B(_05160_),
    .ZN(_01125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10678_ (.A1(\u_cpu.rf_ram.memory[102][7] ),
    .A2(_05150_),
    .ZN(_05161_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10679_ (.A1(_05148_),
    .A2(_05152_),
    .B(_05161_),
    .ZN(_01126_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10680_ (.I(_04958_),
    .Z(_05162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10681_ (.A1(_02876_),
    .A2(_05162_),
    .ZN(_05163_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10682_ (.I(_05163_),
    .Z(_05164_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10683_ (.I(_05163_),
    .Z(_05165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10684_ (.A1(\u_cpu.rf_ram.memory[103][0] ),
    .A2(_05165_),
    .ZN(_05166_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10685_ (.A1(_05130_),
    .A2(_05164_),
    .B(_05166_),
    .ZN(_01127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10686_ (.A1(\u_cpu.rf_ram.memory[103][1] ),
    .A2(_05165_),
    .ZN(_05167_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10687_ (.A1(_05135_),
    .A2(_05164_),
    .B(_05167_),
    .ZN(_01128_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10688_ (.I(_05163_),
    .Z(_05168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10689_ (.A1(\u_cpu.rf_ram.memory[103][2] ),
    .A2(_05168_),
    .ZN(_05169_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10690_ (.A1(_05137_),
    .A2(_05164_),
    .B(_05169_),
    .ZN(_01129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10691_ (.A1(\u_cpu.rf_ram.memory[103][3] ),
    .A2(_05168_),
    .ZN(_05170_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10692_ (.A1(_05140_),
    .A2(_05164_),
    .B(_05170_),
    .ZN(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10693_ (.A1(\u_cpu.rf_ram.memory[103][4] ),
    .A2(_05168_),
    .ZN(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10694_ (.A1(_05142_),
    .A2(_05164_),
    .B(_05171_),
    .ZN(_01131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10695_ (.A1(\u_cpu.rf_ram.memory[103][5] ),
    .A2(_05168_),
    .ZN(_05172_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10696_ (.A1(_05144_),
    .A2(_05165_),
    .B(_05172_),
    .ZN(_01132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10697_ (.A1(\u_cpu.rf_ram.memory[103][6] ),
    .A2(_05168_),
    .ZN(_05173_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10698_ (.A1(_05146_),
    .A2(_05165_),
    .B(_05173_),
    .ZN(_01133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10699_ (.A1(\u_cpu.rf_ram.memory[103][7] ),
    .A2(_05163_),
    .ZN(_05174_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10700_ (.A1(_05148_),
    .A2(_05165_),
    .B(_05174_),
    .ZN(_01134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10701_ (.A1(_03165_),
    .A2(_05162_),
    .ZN(_05175_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10702_ (.I(_05175_),
    .Z(_05176_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10703_ (.I(_05175_),
    .Z(_05177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10704_ (.A1(\u_cpu.rf_ram.memory[104][0] ),
    .A2(_05177_),
    .ZN(_05178_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10705_ (.A1(_05130_),
    .A2(_05176_),
    .B(_05178_),
    .ZN(_01135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10706_ (.A1(\u_cpu.rf_ram.memory[104][1] ),
    .A2(_05177_),
    .ZN(_05179_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10707_ (.A1(_05135_),
    .A2(_05176_),
    .B(_05179_),
    .ZN(_01136_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10708_ (.I(_05175_),
    .Z(_05180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10709_ (.A1(\u_cpu.rf_ram.memory[104][2] ),
    .A2(_05180_),
    .ZN(_05181_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10710_ (.A1(_05137_),
    .A2(_05176_),
    .B(_05181_),
    .ZN(_01137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10711_ (.A1(\u_cpu.rf_ram.memory[104][3] ),
    .A2(_05180_),
    .ZN(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10712_ (.A1(_05140_),
    .A2(_05176_),
    .B(_05182_),
    .ZN(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10713_ (.A1(\u_cpu.rf_ram.memory[104][4] ),
    .A2(_05180_),
    .ZN(_05183_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10714_ (.A1(_05142_),
    .A2(_05176_),
    .B(_05183_),
    .ZN(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10715_ (.A1(\u_cpu.rf_ram.memory[104][5] ),
    .A2(_05180_),
    .ZN(_05184_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10716_ (.A1(_05144_),
    .A2(_05177_),
    .B(_05184_),
    .ZN(_01140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10717_ (.A1(\u_cpu.rf_ram.memory[104][6] ),
    .A2(_05180_),
    .ZN(_05185_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10718_ (.A1(_05146_),
    .A2(_05177_),
    .B(_05185_),
    .ZN(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10719_ (.A1(\u_cpu.rf_ram.memory[104][7] ),
    .A2(_05175_),
    .ZN(_05186_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10720_ (.A1(_05148_),
    .A2(_05177_),
    .B(_05186_),
    .ZN(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10721_ (.A1(_03002_),
    .A2(_05162_),
    .ZN(_05187_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10722_ (.I(_05187_),
    .Z(_05188_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10723_ (.I(_05187_),
    .Z(_05189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10724_ (.A1(\u_cpu.rf_ram.memory[99][0] ),
    .A2(_05189_),
    .ZN(_05190_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10725_ (.A1(_05130_),
    .A2(_05188_),
    .B(_05190_),
    .ZN(_01143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10726_ (.A1(\u_cpu.rf_ram.memory[99][1] ),
    .A2(_05189_),
    .ZN(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10727_ (.A1(_05135_),
    .A2(_05188_),
    .B(_05191_),
    .ZN(_01144_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10728_ (.I(_05187_),
    .Z(_05192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10729_ (.A1(\u_cpu.rf_ram.memory[99][2] ),
    .A2(_05192_),
    .ZN(_05193_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10730_ (.A1(_05137_),
    .A2(_05188_),
    .B(_05193_),
    .ZN(_01145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10731_ (.A1(\u_cpu.rf_ram.memory[99][3] ),
    .A2(_05192_),
    .ZN(_05194_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10732_ (.A1(_05140_),
    .A2(_05188_),
    .B(_05194_),
    .ZN(_01146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10733_ (.A1(\u_cpu.rf_ram.memory[99][4] ),
    .A2(_05192_),
    .ZN(_05195_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10734_ (.A1(_05142_),
    .A2(_05188_),
    .B(_05195_),
    .ZN(_01147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10735_ (.A1(\u_cpu.rf_ram.memory[99][5] ),
    .A2(_05192_),
    .ZN(_05196_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10736_ (.A1(_05144_),
    .A2(_05189_),
    .B(_05196_),
    .ZN(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10737_ (.A1(\u_cpu.rf_ram.memory[99][6] ),
    .A2(_05192_),
    .ZN(_05197_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10738_ (.A1(_05146_),
    .A2(_05189_),
    .B(_05197_),
    .ZN(_01149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10739_ (.A1(\u_cpu.rf_ram.memory[99][7] ),
    .A2(_05187_),
    .ZN(_05198_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10740_ (.A1(_05148_),
    .A2(_05189_),
    .B(_05198_),
    .ZN(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10741_ (.I(_04807_),
    .Z(_05199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10742_ (.A1(_02922_),
    .A2(_03061_),
    .ZN(_05200_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10743_ (.I(_05200_),
    .Z(_05201_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10744_ (.I(_05200_),
    .Z(_05202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10745_ (.A1(\u_cpu.rf_ram.memory[79][0] ),
    .A2(_05202_),
    .ZN(_05203_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10746_ (.A1(_05199_),
    .A2(_05201_),
    .B(_05203_),
    .ZN(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10747_ (.I(_04813_),
    .Z(_05204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10748_ (.A1(\u_cpu.rf_ram.memory[79][1] ),
    .A2(_05202_),
    .ZN(_05205_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10749_ (.A1(_05204_),
    .A2(_05201_),
    .B(_05205_),
    .ZN(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10750_ (.I(_04816_),
    .Z(_05206_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10751_ (.I(_05200_),
    .Z(_05207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10752_ (.A1(\u_cpu.rf_ram.memory[79][2] ),
    .A2(_05207_),
    .ZN(_05208_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10753_ (.A1(_05206_),
    .A2(_05201_),
    .B(_05208_),
    .ZN(_01153_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10754_ (.I(_04820_),
    .Z(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10755_ (.A1(\u_cpu.rf_ram.memory[79][3] ),
    .A2(_05207_),
    .ZN(_05210_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10756_ (.A1(_05209_),
    .A2(_05201_),
    .B(_05210_),
    .ZN(_01154_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10757_ (.I(_04823_),
    .Z(_05211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10758_ (.A1(\u_cpu.rf_ram.memory[79][4] ),
    .A2(_05207_),
    .ZN(_05212_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10759_ (.A1(_05211_),
    .A2(_05201_),
    .B(_05212_),
    .ZN(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10760_ (.I(_04826_),
    .Z(_05213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10761_ (.A1(\u_cpu.rf_ram.memory[79][5] ),
    .A2(_05207_),
    .ZN(_05214_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10762_ (.A1(_05213_),
    .A2(_05202_),
    .B(_05214_),
    .ZN(_01156_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10763_ (.I(_04829_),
    .Z(_05215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10764_ (.A1(\u_cpu.rf_ram.memory[79][6] ),
    .A2(_05207_),
    .ZN(_05216_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10765_ (.A1(_05215_),
    .A2(_05202_),
    .B(_05216_),
    .ZN(_01157_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10766_ (.I(_04832_),
    .Z(_05217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10767_ (.A1(\u_cpu.rf_ram.memory[79][7] ),
    .A2(_05200_),
    .ZN(_05218_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10768_ (.A1(_05217_),
    .A2(_05202_),
    .B(_05218_),
    .ZN(_01158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10769_ (.A1(_03019_),
    .A2(_05162_),
    .ZN(_05219_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10770_ (.I(_05219_),
    .Z(_05220_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10771_ (.I(_05219_),
    .Z(_05221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10772_ (.A1(\u_cpu.rf_ram.memory[105][0] ),
    .A2(_05221_),
    .ZN(_05222_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10773_ (.A1(_05199_),
    .A2(_05220_),
    .B(_05222_),
    .ZN(_01159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10774_ (.A1(\u_cpu.rf_ram.memory[105][1] ),
    .A2(_05221_),
    .ZN(_05223_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10775_ (.A1(_05204_),
    .A2(_05220_),
    .B(_05223_),
    .ZN(_01160_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10776_ (.I(_05219_),
    .Z(_05224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10777_ (.A1(\u_cpu.rf_ram.memory[105][2] ),
    .A2(_05224_),
    .ZN(_05225_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10778_ (.A1(_05206_),
    .A2(_05220_),
    .B(_05225_),
    .ZN(_01161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10779_ (.A1(\u_cpu.rf_ram.memory[105][3] ),
    .A2(_05224_),
    .ZN(_05226_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10780_ (.A1(_05209_),
    .A2(_05220_),
    .B(_05226_),
    .ZN(_01162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10781_ (.A1(\u_cpu.rf_ram.memory[105][4] ),
    .A2(_05224_),
    .ZN(_05227_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10782_ (.A1(_05211_),
    .A2(_05220_),
    .B(_05227_),
    .ZN(_01163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10783_ (.A1(\u_cpu.rf_ram.memory[105][5] ),
    .A2(_05224_),
    .ZN(_05228_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10784_ (.A1(_05213_),
    .A2(_05221_),
    .B(_05228_),
    .ZN(_01164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10785_ (.A1(\u_cpu.rf_ram.memory[105][6] ),
    .A2(_05224_),
    .ZN(_05229_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10786_ (.A1(_05215_),
    .A2(_05221_),
    .B(_05229_),
    .ZN(_01165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10787_ (.A1(\u_cpu.rf_ram.memory[105][7] ),
    .A2(_05219_),
    .ZN(_05230_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10788_ (.A1(_05217_),
    .A2(_05221_),
    .B(_05230_),
    .ZN(_01166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10789_ (.A1(_02937_),
    .A2(_05162_),
    .ZN(_05231_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10790_ (.I(_05231_),
    .Z(_05232_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10791_ (.I(_05231_),
    .Z(_05233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10792_ (.A1(\u_cpu.rf_ram.memory[106][0] ),
    .A2(_05233_),
    .ZN(_05234_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10793_ (.A1(_05199_),
    .A2(_05232_),
    .B(_05234_),
    .ZN(_01167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10794_ (.A1(\u_cpu.rf_ram.memory[106][1] ),
    .A2(_05233_),
    .ZN(_05235_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10795_ (.A1(_05204_),
    .A2(_05232_),
    .B(_05235_),
    .ZN(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10796_ (.I(_05231_),
    .Z(_05236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10797_ (.A1(\u_cpu.rf_ram.memory[106][2] ),
    .A2(_05236_),
    .ZN(_05237_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10798_ (.A1(_05206_),
    .A2(_05232_),
    .B(_05237_),
    .ZN(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10799_ (.A1(\u_cpu.rf_ram.memory[106][3] ),
    .A2(_05236_),
    .ZN(_05238_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10800_ (.A1(_05209_),
    .A2(_05232_),
    .B(_05238_),
    .ZN(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10801_ (.A1(\u_cpu.rf_ram.memory[106][4] ),
    .A2(_05236_),
    .ZN(_05239_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10802_ (.A1(_05211_),
    .A2(_05232_),
    .B(_05239_),
    .ZN(_01171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10803_ (.A1(\u_cpu.rf_ram.memory[106][5] ),
    .A2(_05236_),
    .ZN(_05240_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10804_ (.A1(_05213_),
    .A2(_05233_),
    .B(_05240_),
    .ZN(_01172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10805_ (.A1(\u_cpu.rf_ram.memory[106][6] ),
    .A2(_05236_),
    .ZN(_05241_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10806_ (.A1(_05215_),
    .A2(_05233_),
    .B(_05241_),
    .ZN(_01173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10807_ (.A1(\u_cpu.rf_ram.memory[106][7] ),
    .A2(_05231_),
    .ZN(_05242_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10808_ (.A1(_05217_),
    .A2(_05233_),
    .B(_05242_),
    .ZN(_01174_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10809_ (.I(_04958_),
    .Z(_05243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10810_ (.A1(_03033_),
    .A2(_05243_),
    .ZN(_05244_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10811_ (.I(_05244_),
    .Z(_05245_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10812_ (.I(_05244_),
    .Z(_05246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10813_ (.A1(\u_cpu.rf_ram.memory[107][0] ),
    .A2(_05246_),
    .ZN(_05247_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10814_ (.A1(_05199_),
    .A2(_05245_),
    .B(_05247_),
    .ZN(_01175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10815_ (.A1(\u_cpu.rf_ram.memory[107][1] ),
    .A2(_05246_),
    .ZN(_05248_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10816_ (.A1(_05204_),
    .A2(_05245_),
    .B(_05248_),
    .ZN(_01176_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10817_ (.I(_05244_),
    .Z(_05249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10818_ (.A1(\u_cpu.rf_ram.memory[107][2] ),
    .A2(_05249_),
    .ZN(_05250_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10819_ (.A1(_05206_),
    .A2(_05245_),
    .B(_05250_),
    .ZN(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10820_ (.A1(\u_cpu.rf_ram.memory[107][3] ),
    .A2(_05249_),
    .ZN(_05251_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10821_ (.A1(_05209_),
    .A2(_05245_),
    .B(_05251_),
    .ZN(_01178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10822_ (.A1(\u_cpu.rf_ram.memory[107][4] ),
    .A2(_05249_),
    .ZN(_05252_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10823_ (.A1(_05211_),
    .A2(_05245_),
    .B(_05252_),
    .ZN(_01179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10824_ (.A1(\u_cpu.rf_ram.memory[107][5] ),
    .A2(_05249_),
    .ZN(_05253_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10825_ (.A1(_05213_),
    .A2(_05246_),
    .B(_05253_),
    .ZN(_01180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10826_ (.A1(\u_cpu.rf_ram.memory[107][6] ),
    .A2(_05249_),
    .ZN(_05254_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10827_ (.A1(_05215_),
    .A2(_05246_),
    .B(_05254_),
    .ZN(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10828_ (.A1(\u_cpu.rf_ram.memory[107][7] ),
    .A2(_05244_),
    .ZN(_05255_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10829_ (.A1(_05217_),
    .A2(_05246_),
    .B(_05255_),
    .ZN(_01182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10830_ (.A1(_04091_),
    .A2(_03310_),
    .ZN(_05256_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10831_ (.I(_05256_),
    .Z(_05257_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10832_ (.I(_05256_),
    .Z(_05258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10833_ (.A1(\u_cpu.rf_ram.memory[83][0] ),
    .A2(_05258_),
    .ZN(_05259_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10834_ (.A1(_05199_),
    .A2(_05257_),
    .B(_05259_),
    .ZN(_01183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10835_ (.A1(\u_cpu.rf_ram.memory[83][1] ),
    .A2(_05258_),
    .ZN(_05260_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10836_ (.A1(_05204_),
    .A2(_05257_),
    .B(_05260_),
    .ZN(_01184_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10837_ (.I(_05256_),
    .Z(_05261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10838_ (.A1(\u_cpu.rf_ram.memory[83][2] ),
    .A2(_05261_),
    .ZN(_05262_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10839_ (.A1(_05206_),
    .A2(_05257_),
    .B(_05262_),
    .ZN(_01185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10840_ (.A1(\u_cpu.rf_ram.memory[83][3] ),
    .A2(_05261_),
    .ZN(_05263_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10841_ (.A1(_05209_),
    .A2(_05257_),
    .B(_05263_),
    .ZN(_01186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10842_ (.A1(\u_cpu.rf_ram.memory[83][4] ),
    .A2(_05261_),
    .ZN(_05264_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10843_ (.A1(_05211_),
    .A2(_05257_),
    .B(_05264_),
    .ZN(_01187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10844_ (.A1(\u_cpu.rf_ram.memory[83][5] ),
    .A2(_05261_),
    .ZN(_05265_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10845_ (.A1(_05213_),
    .A2(_05258_),
    .B(_05265_),
    .ZN(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10846_ (.A1(\u_cpu.rf_ram.memory[83][6] ),
    .A2(_05261_),
    .ZN(_05266_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10847_ (.A1(_05215_),
    .A2(_05258_),
    .B(_05266_),
    .ZN(_01189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10848_ (.A1(\u_cpu.rf_ram.memory[83][7] ),
    .A2(_05256_),
    .ZN(_05267_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10849_ (.A1(_05217_),
    .A2(_05258_),
    .B(_05267_),
    .ZN(_01190_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10850_ (.I(_04807_),
    .Z(_05268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10851_ (.A1(_02981_),
    .A2(_05243_),
    .ZN(_05269_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10852_ (.I(_05269_),
    .Z(_05270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10853_ (.I(_05269_),
    .Z(_05271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10854_ (.A1(\u_cpu.rf_ram.memory[108][0] ),
    .A2(_05271_),
    .ZN(_05272_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10855_ (.A1(_05268_),
    .A2(_05270_),
    .B(_05272_),
    .ZN(_01191_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10856_ (.I(_04813_),
    .Z(_05273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10857_ (.A1(\u_cpu.rf_ram.memory[108][1] ),
    .A2(_05271_),
    .ZN(_05274_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10858_ (.A1(_05273_),
    .A2(_05270_),
    .B(_05274_),
    .ZN(_01192_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10859_ (.I(_04816_),
    .Z(_05275_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10860_ (.I(_05269_),
    .Z(_05276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10861_ (.A1(\u_cpu.rf_ram.memory[108][2] ),
    .A2(_05276_),
    .ZN(_05277_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10862_ (.A1(_05275_),
    .A2(_05270_),
    .B(_05277_),
    .ZN(_01193_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10863_ (.I(_04820_),
    .Z(_05278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10864_ (.A1(\u_cpu.rf_ram.memory[108][3] ),
    .A2(_05276_),
    .ZN(_05279_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10865_ (.A1(_05278_),
    .A2(_05270_),
    .B(_05279_),
    .ZN(_01194_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10866_ (.I(_04823_),
    .Z(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10867_ (.A1(\u_cpu.rf_ram.memory[108][4] ),
    .A2(_05276_),
    .ZN(_05281_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10868_ (.A1(_05280_),
    .A2(_05270_),
    .B(_05281_),
    .ZN(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10869_ (.I(_04826_),
    .Z(_05282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10870_ (.A1(\u_cpu.rf_ram.memory[108][5] ),
    .A2(_05276_),
    .ZN(_05283_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10871_ (.A1(_05282_),
    .A2(_05271_),
    .B(_05283_),
    .ZN(_01196_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10872_ (.I(_04829_),
    .Z(_05284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10873_ (.A1(\u_cpu.rf_ram.memory[108][6] ),
    .A2(_05276_),
    .ZN(_05285_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10874_ (.A1(_05284_),
    .A2(_05271_),
    .B(_05285_),
    .ZN(_01197_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10875_ (.I(_04832_),
    .Z(_05286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10876_ (.A1(\u_cpu.rf_ram.memory[108][7] ),
    .A2(_05269_),
    .ZN(_05287_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10877_ (.A1(_05286_),
    .A2(_05271_),
    .B(_05287_),
    .ZN(_01198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10878_ (.A1(_02785_),
    .A2(_03227_),
    .ZN(_05288_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10879_ (.I(_05288_),
    .Z(_05289_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10880_ (.I(_05288_),
    .Z(_05290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10881_ (.A1(\u_cpu.rf_ram.memory[69][0] ),
    .A2(_05290_),
    .ZN(_05291_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10882_ (.A1(_05268_),
    .A2(_05289_),
    .B(_05291_),
    .ZN(_01199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10883_ (.A1(\u_cpu.rf_ram.memory[69][1] ),
    .A2(_05290_),
    .ZN(_05292_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10884_ (.A1(_05273_),
    .A2(_05289_),
    .B(_05292_),
    .ZN(_01200_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10885_ (.I(_05288_),
    .Z(_05293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10886_ (.A1(\u_cpu.rf_ram.memory[69][2] ),
    .A2(_05293_),
    .ZN(_05294_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10887_ (.A1(_05275_),
    .A2(_05289_),
    .B(_05294_),
    .ZN(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10888_ (.A1(\u_cpu.rf_ram.memory[69][3] ),
    .A2(_05293_),
    .ZN(_05295_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10889_ (.A1(_05278_),
    .A2(_05289_),
    .B(_05295_),
    .ZN(_01202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10890_ (.A1(\u_cpu.rf_ram.memory[69][4] ),
    .A2(_05293_),
    .ZN(_05296_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10891_ (.A1(_05280_),
    .A2(_05289_),
    .B(_05296_),
    .ZN(_01203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10892_ (.A1(\u_cpu.rf_ram.memory[69][5] ),
    .A2(_05293_),
    .ZN(_05297_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10893_ (.A1(_05282_),
    .A2(_05290_),
    .B(_05297_),
    .ZN(_01204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10894_ (.A1(\u_cpu.rf_ram.memory[69][6] ),
    .A2(_05293_),
    .ZN(_05298_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10895_ (.A1(_05284_),
    .A2(_05290_),
    .B(_05298_),
    .ZN(_01205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10896_ (.A1(\u_cpu.rf_ram.memory[69][7] ),
    .A2(_05288_),
    .ZN(_05299_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10897_ (.A1(_05286_),
    .A2(_05290_),
    .B(_05299_),
    .ZN(_01206_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10898_ (.I(_02730_),
    .Z(_05300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10899_ (.A1(_05300_),
    .A2(_02831_),
    .ZN(_05301_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10900_ (.I(_05301_),
    .Z(_05302_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10901_ (.I(_05301_),
    .Z(_05303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10902_ (.A1(\u_cpu.rf_ram.memory[84][0] ),
    .A2(_05303_),
    .ZN(_05304_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10903_ (.A1(_05268_),
    .A2(_05302_),
    .B(_05304_),
    .ZN(_01207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10904_ (.A1(\u_cpu.rf_ram.memory[84][1] ),
    .A2(_05303_),
    .ZN(_05305_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10905_ (.A1(_05273_),
    .A2(_05302_),
    .B(_05305_),
    .ZN(_01208_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10906_ (.I(_05301_),
    .Z(_05306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10907_ (.A1(\u_cpu.rf_ram.memory[84][2] ),
    .A2(_05306_),
    .ZN(_05307_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10908_ (.A1(_05275_),
    .A2(_05302_),
    .B(_05307_),
    .ZN(_01209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10909_ (.A1(\u_cpu.rf_ram.memory[84][3] ),
    .A2(_05306_),
    .ZN(_05308_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10910_ (.A1(_05278_),
    .A2(_05302_),
    .B(_05308_),
    .ZN(_01210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10911_ (.A1(\u_cpu.rf_ram.memory[84][4] ),
    .A2(_05306_),
    .ZN(_05309_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10912_ (.A1(_05280_),
    .A2(_05302_),
    .B(_05309_),
    .ZN(_01211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10913_ (.A1(\u_cpu.rf_ram.memory[84][5] ),
    .A2(_05306_),
    .ZN(_05310_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10914_ (.A1(_05282_),
    .A2(_05303_),
    .B(_05310_),
    .ZN(_01212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10915_ (.A1(\u_cpu.rf_ram.memory[84][6] ),
    .A2(_05306_),
    .ZN(_05311_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10916_ (.A1(_05284_),
    .A2(_05303_),
    .B(_05311_),
    .ZN(_01213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10917_ (.A1(\u_cpu.rf_ram.memory[84][7] ),
    .A2(_05301_),
    .ZN(_05312_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10918_ (.A1(_05286_),
    .A2(_05303_),
    .B(_05312_),
    .ZN(_01214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10919_ (.A1(_03004_),
    .A2(_03034_),
    .ZN(_05313_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10920_ (.I(_05313_),
    .Z(_05314_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10921_ (.I(_05313_),
    .Z(_05315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10922_ (.A1(\u_cpu.rf_ram.memory[59][0] ),
    .A2(_05315_),
    .ZN(_05316_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10923_ (.A1(_05268_),
    .A2(_05314_),
    .B(_05316_),
    .ZN(_01215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10924_ (.A1(\u_cpu.rf_ram.memory[59][1] ),
    .A2(_05315_),
    .ZN(_05317_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10925_ (.A1(_05273_),
    .A2(_05314_),
    .B(_05317_),
    .ZN(_01216_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10926_ (.I(_05313_),
    .Z(_05318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10927_ (.A1(\u_cpu.rf_ram.memory[59][2] ),
    .A2(_05318_),
    .ZN(_05319_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10928_ (.A1(_05275_),
    .A2(_05314_),
    .B(_05319_),
    .ZN(_01217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10929_ (.A1(\u_cpu.rf_ram.memory[59][3] ),
    .A2(_05318_),
    .ZN(_05320_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10930_ (.A1(_05278_),
    .A2(_05314_),
    .B(_05320_),
    .ZN(_01218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10931_ (.A1(\u_cpu.rf_ram.memory[59][4] ),
    .A2(_05318_),
    .ZN(_05321_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10932_ (.A1(_05280_),
    .A2(_05314_),
    .B(_05321_),
    .ZN(_01219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10933_ (.A1(\u_cpu.rf_ram.memory[59][5] ),
    .A2(_05318_),
    .ZN(_05322_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10934_ (.A1(_05282_),
    .A2(_05315_),
    .B(_05322_),
    .ZN(_01220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10935_ (.A1(\u_cpu.rf_ram.memory[59][6] ),
    .A2(_05318_),
    .ZN(_05323_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10936_ (.A1(_05284_),
    .A2(_05315_),
    .B(_05323_),
    .ZN(_01221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10937_ (.A1(\u_cpu.rf_ram.memory[59][7] ),
    .A2(_05313_),
    .ZN(_05324_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10938_ (.A1(_05286_),
    .A2(_05315_),
    .B(_05324_),
    .ZN(_01222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10939_ (.A1(_03870_),
    .A2(_02938_),
    .ZN(_05325_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10940_ (.I(_05325_),
    .Z(_05326_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10941_ (.I0(_04184_),
    .I1(\u_cpu.rf_ram.memory[10][0] ),
    .S(_05326_),
    .Z(_05327_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10942_ (.I(_05327_),
    .Z(_01223_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10943_ (.I0(_04188_),
    .I1(\u_cpu.rf_ram.memory[10][1] ),
    .S(_05326_),
    .Z(_05328_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10944_ (.I(_05328_),
    .Z(_01224_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10945_ (.I0(_04190_),
    .I1(\u_cpu.rf_ram.memory[10][2] ),
    .S(_05326_),
    .Z(_05329_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10946_ (.I(_05329_),
    .Z(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10947_ (.I0(_04192_),
    .I1(\u_cpu.rf_ram.memory[10][3] ),
    .S(_05326_),
    .Z(_05330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10948_ (.I(_05330_),
    .Z(_01226_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10949_ (.I0(_04194_),
    .I1(\u_cpu.rf_ram.memory[10][4] ),
    .S(_05326_),
    .Z(_05331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10950_ (.I(_05331_),
    .Z(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10951_ (.I0(_04196_),
    .I1(\u_cpu.rf_ram.memory[10][5] ),
    .S(_05325_),
    .Z(_05332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10952_ (.I(_05332_),
    .Z(_01228_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10953_ (.I0(_04198_),
    .I1(\u_cpu.rf_ram.memory[10][6] ),
    .S(_05325_),
    .Z(_05333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10954_ (.I(_05333_),
    .Z(_01229_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10955_ (.I0(_04200_),
    .I1(\u_cpu.rf_ram.memory[10][7] ),
    .S(_05325_),
    .Z(_05334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10956_ (.I(_05334_),
    .Z(_01230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10957_ (.A1(_05300_),
    .A2(_02786_),
    .ZN(_05335_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10958_ (.I(_05335_),
    .Z(_05336_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10959_ (.I(_05335_),
    .Z(_05337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10960_ (.A1(\u_cpu.rf_ram.memory[85][0] ),
    .A2(_05337_),
    .ZN(_05338_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10961_ (.A1(_05268_),
    .A2(_05336_),
    .B(_05338_),
    .ZN(_01231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10962_ (.A1(\u_cpu.rf_ram.memory[85][1] ),
    .A2(_05337_),
    .ZN(_05339_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10963_ (.A1(_05273_),
    .A2(_05336_),
    .B(_05339_),
    .ZN(_01232_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10964_ (.I(_05335_),
    .Z(_05340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10965_ (.A1(\u_cpu.rf_ram.memory[85][2] ),
    .A2(_05340_),
    .ZN(_05341_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10966_ (.A1(_05275_),
    .A2(_05336_),
    .B(_05341_),
    .ZN(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10967_ (.A1(\u_cpu.rf_ram.memory[85][3] ),
    .A2(_05340_),
    .ZN(_05342_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10968_ (.A1(_05278_),
    .A2(_05336_),
    .B(_05342_),
    .ZN(_01234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10969_ (.A1(\u_cpu.rf_ram.memory[85][4] ),
    .A2(_05340_),
    .ZN(_05343_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10970_ (.A1(_05280_),
    .A2(_05336_),
    .B(_05343_),
    .ZN(_01235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10971_ (.A1(\u_cpu.rf_ram.memory[85][5] ),
    .A2(_05340_),
    .ZN(_05344_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10972_ (.A1(_05282_),
    .A2(_05337_),
    .B(_05344_),
    .ZN(_01236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10973_ (.A1(\u_cpu.rf_ram.memory[85][6] ),
    .A2(_05340_),
    .ZN(_05345_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10974_ (.A1(_05284_),
    .A2(_05337_),
    .B(_05345_),
    .ZN(_01237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10975_ (.A1(\u_cpu.rf_ram.memory[85][7] ),
    .A2(_05335_),
    .ZN(_05346_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10976_ (.A1(_05286_),
    .A2(_05337_),
    .B(_05346_),
    .ZN(_01238_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10977_ (.I(_02739_),
    .Z(_05347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10978_ (.A1(_02920_),
    .A2(_05243_),
    .ZN(_05348_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10979_ (.I(_05348_),
    .Z(_05349_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10980_ (.I(_05348_),
    .Z(_05350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10981_ (.A1(\u_cpu.rf_ram.memory[110][0] ),
    .A2(_05350_),
    .ZN(_05351_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10982_ (.A1(_05347_),
    .A2(_05349_),
    .B(_05351_),
    .ZN(_01239_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10983_ (.I(_02745_),
    .Z(_05352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10984_ (.A1(\u_cpu.rf_ram.memory[110][1] ),
    .A2(_05350_),
    .ZN(_05353_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10985_ (.A1(_05352_),
    .A2(_05349_),
    .B(_05353_),
    .ZN(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10986_ (.I(_02751_),
    .Z(_05354_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10987_ (.I(_05348_),
    .Z(_05355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10988_ (.A1(\u_cpu.rf_ram.memory[110][2] ),
    .A2(_05355_),
    .ZN(_05356_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10989_ (.A1(_05354_),
    .A2(_05349_),
    .B(_05356_),
    .ZN(_01241_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10990_ (.I(_02757_),
    .Z(_05357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10991_ (.A1(\u_cpu.rf_ram.memory[110][3] ),
    .A2(_05355_),
    .ZN(_05358_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10992_ (.A1(_05357_),
    .A2(_05349_),
    .B(_05358_),
    .ZN(_01242_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10993_ (.I(_02762_),
    .Z(_05359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10994_ (.A1(\u_cpu.rf_ram.memory[110][4] ),
    .A2(_05355_),
    .ZN(_05360_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10995_ (.A1(_05359_),
    .A2(_05349_),
    .B(_05360_),
    .ZN(_01243_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10996_ (.I(_02767_),
    .Z(_05361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10997_ (.A1(\u_cpu.rf_ram.memory[110][5] ),
    .A2(_05355_),
    .ZN(_05362_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10998_ (.A1(_05361_),
    .A2(_05350_),
    .B(_05362_),
    .ZN(_01244_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10999_ (.I(_02772_),
    .Z(_05363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11000_ (.A1(\u_cpu.rf_ram.memory[110][6] ),
    .A2(_05355_),
    .ZN(_05364_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11001_ (.A1(_05363_),
    .A2(_05350_),
    .B(_05364_),
    .ZN(_01245_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11002_ (.I(_02777_),
    .Z(_05365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11003_ (.A1(\u_cpu.rf_ram.memory[110][7] ),
    .A2(_05348_),
    .ZN(_05366_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11004_ (.A1(_05365_),
    .A2(_05350_),
    .B(_05366_),
    .ZN(_01246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11005_ (.A1(_05300_),
    .A2(_03286_),
    .ZN(_05367_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11006_ (.I(_05367_),
    .Z(_05368_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11007_ (.I(_05367_),
    .Z(_05369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11008_ (.A1(\u_cpu.rf_ram.memory[86][0] ),
    .A2(_05369_),
    .ZN(_05370_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11009_ (.A1(_05347_),
    .A2(_05368_),
    .B(_05370_),
    .ZN(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11010_ (.A1(\u_cpu.rf_ram.memory[86][1] ),
    .A2(_05369_),
    .ZN(_05371_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11011_ (.A1(_05352_),
    .A2(_05368_),
    .B(_05371_),
    .ZN(_01248_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11012_ (.I(_05367_),
    .Z(_05372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11013_ (.A1(\u_cpu.rf_ram.memory[86][2] ),
    .A2(_05372_),
    .ZN(_05373_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11014_ (.A1(_05354_),
    .A2(_05368_),
    .B(_05373_),
    .ZN(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11015_ (.A1(\u_cpu.rf_ram.memory[86][3] ),
    .A2(_05372_),
    .ZN(_05374_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11016_ (.A1(_05357_),
    .A2(_05368_),
    .B(_05374_),
    .ZN(_01250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11017_ (.A1(\u_cpu.rf_ram.memory[86][4] ),
    .A2(_05372_),
    .ZN(_05375_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11018_ (.A1(_05359_),
    .A2(_05368_),
    .B(_05375_),
    .ZN(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11019_ (.A1(\u_cpu.rf_ram.memory[86][5] ),
    .A2(_05372_),
    .ZN(_05376_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11020_ (.A1(_05361_),
    .A2(_05369_),
    .B(_05376_),
    .ZN(_01252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11021_ (.A1(\u_cpu.rf_ram.memory[86][6] ),
    .A2(_05372_),
    .ZN(_05377_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11022_ (.A1(_05363_),
    .A2(_05369_),
    .B(_05377_),
    .ZN(_01253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11023_ (.A1(\u_cpu.rf_ram.memory[86][7] ),
    .A2(_05367_),
    .ZN(_05378_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11024_ (.A1(_05365_),
    .A2(_05369_),
    .B(_05378_),
    .ZN(_01254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11025_ (.A1(_03061_),
    .A2(_05243_),
    .ZN(_05379_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11026_ (.I(_05379_),
    .Z(_05380_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11027_ (.I(_05379_),
    .Z(_05381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11028_ (.A1(\u_cpu.rf_ram.memory[111][0] ),
    .A2(_05381_),
    .ZN(_05382_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11029_ (.A1(_05347_),
    .A2(_05380_),
    .B(_05382_),
    .ZN(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11030_ (.A1(\u_cpu.rf_ram.memory[111][1] ),
    .A2(_05381_),
    .ZN(_05383_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11031_ (.A1(_05352_),
    .A2(_05380_),
    .B(_05383_),
    .ZN(_01256_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11032_ (.I(_05379_),
    .Z(_05384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11033_ (.A1(\u_cpu.rf_ram.memory[111][2] ),
    .A2(_05384_),
    .ZN(_05385_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11034_ (.A1(_05354_),
    .A2(_05380_),
    .B(_05385_),
    .ZN(_01257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11035_ (.A1(\u_cpu.rf_ram.memory[111][3] ),
    .A2(_05384_),
    .ZN(_05386_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11036_ (.A1(_05357_),
    .A2(_05380_),
    .B(_05386_),
    .ZN(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11037_ (.A1(\u_cpu.rf_ram.memory[111][4] ),
    .A2(_05384_),
    .ZN(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11038_ (.A1(_05359_),
    .A2(_05380_),
    .B(_05387_),
    .ZN(_01259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11039_ (.A1(\u_cpu.rf_ram.memory[111][5] ),
    .A2(_05384_),
    .ZN(_05388_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11040_ (.A1(_05361_),
    .A2(_05381_),
    .B(_05388_),
    .ZN(_01260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11041_ (.A1(\u_cpu.rf_ram.memory[111][6] ),
    .A2(_05384_),
    .ZN(_05389_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11042_ (.A1(_05363_),
    .A2(_05381_),
    .B(_05389_),
    .ZN(_01261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11043_ (.A1(\u_cpu.rf_ram.memory[111][7] ),
    .A2(_05379_),
    .ZN(_05390_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11044_ (.A1(_05365_),
    .A2(_05381_),
    .B(_05390_),
    .ZN(_01262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11045_ (.A1(_05300_),
    .A2(_02877_),
    .ZN(_05391_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11046_ (.I(_05391_),
    .Z(_05392_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11047_ (.I(_05391_),
    .Z(_05393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11048_ (.A1(\u_cpu.rf_ram.memory[87][0] ),
    .A2(_05393_),
    .ZN(_05394_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11049_ (.A1(_05347_),
    .A2(_05392_),
    .B(_05394_),
    .ZN(_01263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11050_ (.A1(\u_cpu.rf_ram.memory[87][1] ),
    .A2(_05393_),
    .ZN(_05395_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11051_ (.A1(_05352_),
    .A2(_05392_),
    .B(_05395_),
    .ZN(_01264_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11052_ (.I(_05391_),
    .Z(_05396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11053_ (.A1(\u_cpu.rf_ram.memory[87][2] ),
    .A2(_05396_),
    .ZN(_05397_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11054_ (.A1(_05354_),
    .A2(_05392_),
    .B(_05397_),
    .ZN(_01265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11055_ (.A1(\u_cpu.rf_ram.memory[87][3] ),
    .A2(_05396_),
    .ZN(_05398_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11056_ (.A1(_05357_),
    .A2(_05392_),
    .B(_05398_),
    .ZN(_01266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11057_ (.A1(\u_cpu.rf_ram.memory[87][4] ),
    .A2(_05396_),
    .ZN(_05399_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11058_ (.A1(_05359_),
    .A2(_05392_),
    .B(_05399_),
    .ZN(_01267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11059_ (.A1(\u_cpu.rf_ram.memory[87][5] ),
    .A2(_05396_),
    .ZN(_05400_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11060_ (.A1(_05361_),
    .A2(_05393_),
    .B(_05400_),
    .ZN(_01268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11061_ (.A1(\u_cpu.rf_ram.memory[87][6] ),
    .A2(_05396_),
    .ZN(_05401_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11062_ (.A1(_05363_),
    .A2(_05393_),
    .B(_05401_),
    .ZN(_01269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11063_ (.A1(\u_cpu.rf_ram.memory[87][7] ),
    .A2(_05391_),
    .ZN(_05402_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11064_ (.A1(_05365_),
    .A2(_05393_),
    .B(_05402_),
    .ZN(_01270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11065_ (.A1(_05300_),
    .A2(_03166_),
    .ZN(_05403_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11066_ (.I(_05403_),
    .Z(_05404_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11067_ (.I(_05403_),
    .Z(_05405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11068_ (.A1(\u_cpu.rf_ram.memory[88][0] ),
    .A2(_05405_),
    .ZN(_05406_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11069_ (.A1(_05347_),
    .A2(_05404_),
    .B(_05406_),
    .ZN(_01271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11070_ (.A1(\u_cpu.rf_ram.memory[88][1] ),
    .A2(_05405_),
    .ZN(_05407_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11071_ (.A1(_05352_),
    .A2(_05404_),
    .B(_05407_),
    .ZN(_01272_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11072_ (.I(_05403_),
    .Z(_05408_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11073_ (.A1(\u_cpu.rf_ram.memory[88][2] ),
    .A2(_05408_),
    .ZN(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11074_ (.A1(_05354_),
    .A2(_05404_),
    .B(_05409_),
    .ZN(_01273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11075_ (.A1(\u_cpu.rf_ram.memory[88][3] ),
    .A2(_05408_),
    .ZN(_05410_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11076_ (.A1(_05357_),
    .A2(_05404_),
    .B(_05410_),
    .ZN(_01274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11077_ (.A1(\u_cpu.rf_ram.memory[88][4] ),
    .A2(_05408_),
    .ZN(_05411_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11078_ (.A1(_05359_),
    .A2(_05404_),
    .B(_05411_),
    .ZN(_01275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11079_ (.A1(\u_cpu.rf_ram.memory[88][5] ),
    .A2(_05408_),
    .ZN(_05412_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11080_ (.A1(_05361_),
    .A2(_05405_),
    .B(_05412_),
    .ZN(_01276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11081_ (.A1(\u_cpu.rf_ram.memory[88][6] ),
    .A2(_05408_),
    .ZN(_05413_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11082_ (.A1(_05363_),
    .A2(_05405_),
    .B(_05413_),
    .ZN(_01277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11083_ (.A1(\u_cpu.rf_ram.memory[88][7] ),
    .A2(_05403_),
    .ZN(_05414_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11084_ (.A1(_05365_),
    .A2(_05405_),
    .B(_05414_),
    .ZN(_01278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11085_ (.A1(_04026_),
    .A2(_02579_),
    .ZN(_05415_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11086_ (.A1(_02529_),
    .A2(_02572_),
    .A3(_02565_),
    .ZN(_05416_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11087_ (.A1(_05415_),
    .A2(_05416_),
    .Z(_05417_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11088_ (.I(_05417_),
    .Z(_05418_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11089_ (.A1(_02693_),
    .A2(_01393_),
    .ZN(_05419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11090_ (.A1(_01386_),
    .A2(\u_cpu.cpu.genblk3.csr.mcause3_0[1] ),
    .ZN(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11091_ (.A1(_05419_),
    .A2(_05420_),
    .ZN(_05421_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11092_ (.A1(_05418_),
    .A2(_05421_),
    .ZN(_05422_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11093_ (.A1(_02568_),
    .A2(_05418_),
    .B(_05422_),
    .ZN(_01279_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11094_ (.A1(_02684_),
    .A2(_02633_),
    .B1(\u_cpu.cpu.genblk3.csr.mcause3_0[2] ),
    .B2(_01386_),
    .ZN(_05423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11095_ (.A1(_05419_),
    .A2(_05423_),
    .ZN(_05424_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11096_ (.I0(_05424_),
    .I1(\u_cpu.cpu.genblk3.csr.mcause3_0[1] ),
    .S(_05417_),
    .Z(_05425_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11097_ (.I(_05425_),
    .Z(_01280_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11098_ (.A1(\u_cpu.cpu.genblk3.csr.mcause3_0[3] ),
    .A2(_01394_),
    .B(_02693_),
    .C(_02684_),
    .ZN(_05426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11099_ (.A1(\u_cpu.cpu.genblk3.csr.mcause3_0[2] ),
    .A2(_05418_),
    .ZN(_05427_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11100_ (.A1(_05418_),
    .A2(_05426_),
    .B(_05427_),
    .ZN(_01281_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11101_ (.I(\u_cpu.cpu.genblk3.csr.mcause3_0[3] ),
    .ZN(_05428_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11102_ (.A1(_01382_),
    .A2(_01393_),
    .B(_05417_),
    .ZN(_05429_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11103_ (.A1(_05428_),
    .A2(_05418_),
    .B1(_05429_),
    .B2(_02577_),
    .ZN(_01282_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11104_ (.I(\u_cpu.cpu.genblk3.csr.mcause31 ),
    .ZN(_05430_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11105_ (.A1(_04026_),
    .A2(_02572_),
    .B(_02579_),
    .ZN(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11106_ (.A1(_02693_),
    .A2(_05431_),
    .ZN(_05432_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11107_ (.A1(_05430_),
    .A2(_05431_),
    .B1(_05432_),
    .B2(_02577_),
    .ZN(_01283_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11108_ (.I0(\u_cpu.cpu.genblk3.csr.mstatus_mie ),
    .I1(\u_cpu.cpu.genblk3.csr.mstatus_mpie ),
    .S(_05415_),
    .Z(_05433_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11109_ (.I(_05433_),
    .Z(_01284_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11110_ (.I(\u_cpu.cpu.genblk3.csr.mie_mtie ),
    .ZN(_05434_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _11111_ (.A1(\u_cpu.cpu.decode.co_ebreak ),
    .A2(_04034_),
    .A3(_04031_),
    .A4(_02562_),
    .ZN(_05435_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11112_ (.A1(_02566_),
    .A2(_04030_),
    .A3(_05435_),
    .ZN(_05436_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11113_ (.A1(_02576_),
    .A2(_05436_),
    .B(_04032_),
    .ZN(_05437_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11114_ (.A1(_05434_),
    .A2(_05436_),
    .B(_05437_),
    .ZN(_01285_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11115_ (.A1(_04952_),
    .A2(_02576_),
    .ZN(_05438_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11116_ (.A1(\u_cpu.cpu.genblk3.csr.mstatus_mpie ),
    .A2(_01378_),
    .B(_01394_),
    .ZN(_05439_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11117_ (.A1(_04952_),
    .A2(_02567_),
    .ZN(_05440_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11118_ (.A1(\u_cpu.cpu.genblk3.csr.mstatus_mie ),
    .A2(_05415_),
    .A3(_05440_),
    .ZN(_05441_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _11119_ (.A1(_05438_),
    .A2(_05439_),
    .A3(_05440_),
    .B(_05441_),
    .ZN(_01286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11120_ (.A1(\u_cpu.cpu.ctrl.i_iscomp ),
    .A2(_04467_),
    .ZN(_05442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11121_ (.A1(_04494_),
    .A2(_05442_),
    .ZN(_01287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11122_ (.A1(_02693_),
    .A2(_04038_),
    .ZN(_05443_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _11123_ (.A1(_03111_),
    .A2(\u_cpu.cpu.genblk3.csr.timer_irq_r ),
    .A3(_04806_),
    .B(_05443_),
    .ZN(_01288_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11124_ (.I(_02739_),
    .Z(_05444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11125_ (.A1(_05098_),
    .A2(_03033_),
    .ZN(_05445_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11126_ (.I(_05445_),
    .Z(_05446_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11127_ (.I(_05445_),
    .Z(_05447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11128_ (.A1(\u_cpu.rf_ram.memory[27][0] ),
    .A2(_05447_),
    .ZN(_05448_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11129_ (.A1(_05444_),
    .A2(_05446_),
    .B(_05448_),
    .ZN(_01289_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11130_ (.I(_02745_),
    .Z(_05449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11131_ (.A1(\u_cpu.rf_ram.memory[27][1] ),
    .A2(_05447_),
    .ZN(_05450_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11132_ (.A1(_05449_),
    .A2(_05446_),
    .B(_05450_),
    .ZN(_01290_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11133_ (.I(_02751_),
    .Z(_05451_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11134_ (.I(_05445_),
    .Z(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11135_ (.A1(\u_cpu.rf_ram.memory[27][2] ),
    .A2(_05452_),
    .ZN(_05453_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11136_ (.A1(_05451_),
    .A2(_05446_),
    .B(_05453_),
    .ZN(_01291_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11137_ (.I(_02757_),
    .Z(_05454_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11138_ (.A1(\u_cpu.rf_ram.memory[27][3] ),
    .A2(_05452_),
    .ZN(_05455_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11139_ (.A1(_05454_),
    .A2(_05446_),
    .B(_05455_),
    .ZN(_01292_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11140_ (.I(_02762_),
    .Z(_05456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11141_ (.A1(\u_cpu.rf_ram.memory[27][4] ),
    .A2(_05452_),
    .ZN(_05457_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11142_ (.A1(_05456_),
    .A2(_05446_),
    .B(_05457_),
    .ZN(_01293_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11143_ (.I(_02767_),
    .Z(_05458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11144_ (.A1(\u_cpu.rf_ram.memory[27][5] ),
    .A2(_05452_),
    .ZN(_05459_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11145_ (.A1(_05458_),
    .A2(_05447_),
    .B(_05459_),
    .ZN(_01294_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11146_ (.I(_02772_),
    .Z(_05460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11147_ (.A1(\u_cpu.rf_ram.memory[27][6] ),
    .A2(_05452_),
    .ZN(_05461_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11148_ (.A1(_05460_),
    .A2(_05447_),
    .B(_05461_),
    .ZN(_01295_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11149_ (.I(_02777_),
    .Z(_05462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11150_ (.A1(\u_cpu.rf_ram.memory[27][7] ),
    .A2(_05445_),
    .ZN(_05463_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11151_ (.A1(_05462_),
    .A2(_05447_),
    .B(_05463_),
    .ZN(_01296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11152_ (.A1(_05098_),
    .A2(_02938_),
    .ZN(_05464_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11153_ (.I(_05464_),
    .Z(_05465_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11154_ (.I(_05464_),
    .Z(_05466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11155_ (.A1(\u_cpu.rf_ram.memory[26][0] ),
    .A2(_05466_),
    .ZN(_05467_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11156_ (.A1(_05444_),
    .A2(_05465_),
    .B(_05467_),
    .ZN(_01297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11157_ (.A1(\u_cpu.rf_ram.memory[26][1] ),
    .A2(_05466_),
    .ZN(_05468_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11158_ (.A1(_05449_),
    .A2(_05465_),
    .B(_05468_),
    .ZN(_01298_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11159_ (.I(_05464_),
    .Z(_05469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11160_ (.A1(\u_cpu.rf_ram.memory[26][2] ),
    .A2(_05469_),
    .ZN(_05470_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11161_ (.A1(_05451_),
    .A2(_05465_),
    .B(_05470_),
    .ZN(_01299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11162_ (.A1(\u_cpu.rf_ram.memory[26][3] ),
    .A2(_05469_),
    .ZN(_05471_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11163_ (.A1(_05454_),
    .A2(_05465_),
    .B(_05471_),
    .ZN(_01300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11164_ (.A1(\u_cpu.rf_ram.memory[26][4] ),
    .A2(_05469_),
    .ZN(_05472_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11165_ (.A1(_05456_),
    .A2(_05465_),
    .B(_05472_),
    .ZN(_01301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11166_ (.A1(\u_cpu.rf_ram.memory[26][5] ),
    .A2(_05469_),
    .ZN(_05473_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11167_ (.A1(_05458_),
    .A2(_05466_),
    .B(_05473_),
    .ZN(_01302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11168_ (.A1(\u_cpu.rf_ram.memory[26][6] ),
    .A2(_05469_),
    .ZN(_05474_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11169_ (.A1(_05460_),
    .A2(_05466_),
    .B(_05474_),
    .ZN(_01303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11170_ (.A1(\u_cpu.rf_ram.memory[26][7] ),
    .A2(_05464_),
    .ZN(_05475_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11171_ (.A1(_05462_),
    .A2(_05466_),
    .B(_05475_),
    .ZN(_01304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11172_ (.A1(_05098_),
    .A2(_03020_),
    .ZN(_05476_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11173_ (.I(_05476_),
    .Z(_05477_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11174_ (.I(_05476_),
    .Z(_05478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11175_ (.A1(\u_cpu.rf_ram.memory[25][0] ),
    .A2(_05478_),
    .ZN(_05479_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11176_ (.A1(_05444_),
    .A2(_05477_),
    .B(_05479_),
    .ZN(_01305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11177_ (.A1(\u_cpu.rf_ram.memory[25][1] ),
    .A2(_05478_),
    .ZN(_05480_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11178_ (.A1(_05449_),
    .A2(_05477_),
    .B(_05480_),
    .ZN(_01306_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11179_ (.I(_05476_),
    .Z(_05481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11180_ (.A1(\u_cpu.rf_ram.memory[25][2] ),
    .A2(_05481_),
    .ZN(_05482_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11181_ (.A1(_05451_),
    .A2(_05477_),
    .B(_05482_),
    .ZN(_01307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11182_ (.A1(\u_cpu.rf_ram.memory[25][3] ),
    .A2(_05481_),
    .ZN(_05483_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11183_ (.A1(_05454_),
    .A2(_05477_),
    .B(_05483_),
    .ZN(_01308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11184_ (.A1(\u_cpu.rf_ram.memory[25][4] ),
    .A2(_05481_),
    .ZN(_05484_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11185_ (.A1(_05456_),
    .A2(_05477_),
    .B(_05484_),
    .ZN(_01309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11186_ (.A1(\u_cpu.rf_ram.memory[25][5] ),
    .A2(_05481_),
    .ZN(_05485_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11187_ (.A1(_05458_),
    .A2(_05478_),
    .B(_05485_),
    .ZN(_01310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11188_ (.A1(\u_cpu.rf_ram.memory[25][6] ),
    .A2(_05481_),
    .ZN(_05486_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11189_ (.A1(_05460_),
    .A2(_05478_),
    .B(_05486_),
    .ZN(_01311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11190_ (.A1(\u_cpu.rf_ram.memory[25][7] ),
    .A2(_05476_),
    .ZN(_05487_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11191_ (.A1(_05462_),
    .A2(_05478_),
    .B(_05487_),
    .ZN(_01312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11192_ (.A1(_05098_),
    .A2(_03165_),
    .ZN(_05488_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11193_ (.I(_05488_),
    .Z(_05489_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11194_ (.I(_05488_),
    .Z(_05490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11195_ (.A1(\u_cpu.rf_ram.memory[24][0] ),
    .A2(_05490_),
    .ZN(_05491_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11196_ (.A1(_05444_),
    .A2(_05489_),
    .B(_05491_),
    .ZN(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11197_ (.A1(\u_cpu.rf_ram.memory[24][1] ),
    .A2(_05490_),
    .ZN(_05492_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11198_ (.A1(_05449_),
    .A2(_05489_),
    .B(_05492_),
    .ZN(_01314_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11199_ (.I(_05488_),
    .Z(_05493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11200_ (.A1(\u_cpu.rf_ram.memory[24][2] ),
    .A2(_05493_),
    .ZN(_05494_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11201_ (.A1(_05451_),
    .A2(_05489_),
    .B(_05494_),
    .ZN(_01315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11202_ (.A1(\u_cpu.rf_ram.memory[24][3] ),
    .A2(_05493_),
    .ZN(_05495_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11203_ (.A1(_05454_),
    .A2(_05489_),
    .B(_05495_),
    .ZN(_01316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11204_ (.A1(\u_cpu.rf_ram.memory[24][4] ),
    .A2(_05493_),
    .ZN(_05496_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11205_ (.A1(_05456_),
    .A2(_05489_),
    .B(_05496_),
    .ZN(_01317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11206_ (.A1(\u_cpu.rf_ram.memory[24][5] ),
    .A2(_05493_),
    .ZN(_05497_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11207_ (.A1(_05458_),
    .A2(_05490_),
    .B(_05497_),
    .ZN(_01318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11208_ (.A1(\u_cpu.rf_ram.memory[24][6] ),
    .A2(_05493_),
    .ZN(_05498_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11209_ (.A1(_05460_),
    .A2(_05490_),
    .B(_05498_),
    .ZN(_01319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11210_ (.A1(\u_cpu.rf_ram.memory[24][7] ),
    .A2(_05488_),
    .ZN(_05499_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11211_ (.A1(_05462_),
    .A2(_05490_),
    .B(_05499_),
    .ZN(_01320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11212_ (.A1(_02849_),
    .A2(_02891_),
    .ZN(_05500_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11213_ (.I(_05500_),
    .Z(_05501_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11214_ (.I0(_02845_),
    .I1(\u_cpu.rf_ram.memory[0][0] ),
    .S(_05501_),
    .Z(_05502_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11215_ (.I(_05502_),
    .Z(_01321_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11216_ (.I0(_02854_),
    .I1(\u_cpu.rf_ram.memory[0][1] ),
    .S(_05501_),
    .Z(_05503_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11217_ (.I(_05503_),
    .Z(_01322_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11218_ (.I0(_02857_),
    .I1(\u_cpu.rf_ram.memory[0][2] ),
    .S(_05501_),
    .Z(_05504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11219_ (.I(_05504_),
    .Z(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11220_ (.I0(_02860_),
    .I1(\u_cpu.rf_ram.memory[0][3] ),
    .S(_05501_),
    .Z(_05505_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11221_ (.I(_05505_),
    .Z(_01324_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11222_ (.I0(_02863_),
    .I1(\u_cpu.rf_ram.memory[0][4] ),
    .S(_05501_),
    .Z(_05506_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11223_ (.I(_05506_),
    .Z(_01325_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11224_ (.I0(_02866_),
    .I1(\u_cpu.rf_ram.memory[0][5] ),
    .S(_05500_),
    .Z(_05507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11225_ (.I(_05507_),
    .Z(_01326_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11226_ (.I0(_02869_),
    .I1(\u_cpu.rf_ram.memory[0][6] ),
    .S(_05500_),
    .Z(_05508_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11227_ (.I(_05508_),
    .Z(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11228_ (.I0(_02872_),
    .I1(\u_cpu.rf_ram.memory[0][7] ),
    .S(_05500_),
    .Z(_05509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11229_ (.I(_05509_),
    .Z(_01328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11230_ (.A1(_02722_),
    .A2(_05243_),
    .ZN(_05510_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11231_ (.I(_05510_),
    .Z(_05511_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11232_ (.I(_05510_),
    .Z(_05512_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11233_ (.A1(\u_cpu.rf_ram.memory[98][0] ),
    .A2(_05512_),
    .ZN(_05513_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11234_ (.A1(_05444_),
    .A2(_05511_),
    .B(_05513_),
    .ZN(_01329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11235_ (.A1(\u_cpu.rf_ram.memory[98][1] ),
    .A2(_05512_),
    .ZN(_05514_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11236_ (.A1(_05449_),
    .A2(_05511_),
    .B(_05514_),
    .ZN(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11237_ (.I(_05510_),
    .Z(_05515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11238_ (.A1(\u_cpu.rf_ram.memory[98][2] ),
    .A2(_05515_),
    .ZN(_05516_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11239_ (.A1(_05451_),
    .A2(_05511_),
    .B(_05516_),
    .ZN(_01331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11240_ (.A1(\u_cpu.rf_ram.memory[98][3] ),
    .A2(_05515_),
    .ZN(_05517_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11241_ (.A1(_05454_),
    .A2(_05511_),
    .B(_05517_),
    .ZN(_01332_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11242_ (.A1(\u_cpu.rf_ram.memory[98][4] ),
    .A2(_05515_),
    .ZN(_05518_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11243_ (.A1(_05456_),
    .A2(_05511_),
    .B(_05518_),
    .ZN(_01333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11244_ (.A1(\u_cpu.rf_ram.memory[98][5] ),
    .A2(_05515_),
    .ZN(_05519_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11245_ (.A1(_05458_),
    .A2(_05512_),
    .B(_05519_),
    .ZN(_01334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11246_ (.A1(\u_cpu.rf_ram.memory[98][6] ),
    .A2(_05515_),
    .ZN(_05520_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11247_ (.A1(_05460_),
    .A2(_05512_),
    .B(_05520_),
    .ZN(_01335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11248_ (.A1(\u_cpu.rf_ram.memory[98][7] ),
    .A2(_05510_),
    .ZN(_05521_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11249_ (.A1(_05462_),
    .A2(_05512_),
    .B(_05521_),
    .ZN(_01336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11250_ (.A1(_02830_),
    .A2(_04958_),
    .ZN(_05522_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11251_ (.I(_05522_),
    .Z(_05523_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11252_ (.I(_05522_),
    .Z(_05524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11253_ (.A1(\u_cpu.rf_ram.memory[100][0] ),
    .A2(_05524_),
    .ZN(_05525_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11254_ (.A1(_02888_),
    .A2(_05523_),
    .B(_05525_),
    .ZN(_01337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11255_ (.A1(\u_cpu.rf_ram.memory[100][1] ),
    .A2(_05524_),
    .ZN(_05526_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11256_ (.A1(_02896_),
    .A2(_05523_),
    .B(_05526_),
    .ZN(_01338_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11257_ (.I(_05522_),
    .Z(_05527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11258_ (.A1(\u_cpu.rf_ram.memory[100][2] ),
    .A2(_05527_),
    .ZN(_05528_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11259_ (.A1(_02899_),
    .A2(_05523_),
    .B(_05528_),
    .ZN(_01339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11260_ (.A1(\u_cpu.rf_ram.memory[100][3] ),
    .A2(_05527_),
    .ZN(_05529_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11261_ (.A1(_02903_),
    .A2(_05523_),
    .B(_05529_),
    .ZN(_01340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11262_ (.A1(\u_cpu.rf_ram.memory[100][4] ),
    .A2(_05527_),
    .ZN(_05530_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11263_ (.A1(_02906_),
    .A2(_05523_),
    .B(_05530_),
    .ZN(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11264_ (.A1(\u_cpu.rf_ram.memory[100][5] ),
    .A2(_05527_),
    .ZN(_05531_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11265_ (.A1(_02909_),
    .A2(_05524_),
    .B(_05531_),
    .ZN(_01342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11266_ (.A1(\u_cpu.rf_ram.memory[100][6] ),
    .A2(_05527_),
    .ZN(_05532_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11267_ (.A1(_02912_),
    .A2(_05524_),
    .B(_05532_),
    .ZN(_01343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11268_ (.A1(\u_cpu.rf_ram.memory[100][7] ),
    .A2(_05522_),
    .ZN(_05533_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11269_ (.A1(_02915_),
    .A2(_05524_),
    .B(_05533_),
    .ZN(_01344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11270_ (.A1(_02730_),
    .A2(_03019_),
    .ZN(_05534_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11271_ (.I(_05534_),
    .Z(_05535_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11272_ (.I(_05534_),
    .Z(_05536_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11273_ (.A1(\u_cpu.rf_ram.memory[89][0] ),
    .A2(_05536_),
    .ZN(_05537_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11274_ (.A1(_02888_),
    .A2(_05535_),
    .B(_05537_),
    .ZN(_01345_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11275_ (.A1(\u_cpu.rf_ram.memory[89][1] ),
    .A2(_05536_),
    .ZN(_05538_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11276_ (.A1(_02896_),
    .A2(_05535_),
    .B(_05538_),
    .ZN(_01346_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11277_ (.I(_05534_),
    .Z(_05539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11278_ (.A1(\u_cpu.rf_ram.memory[89][2] ),
    .A2(_05539_),
    .ZN(_05540_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11279_ (.A1(_02899_),
    .A2(_05535_),
    .B(_05540_),
    .ZN(_01347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11280_ (.A1(\u_cpu.rf_ram.memory[89][3] ),
    .A2(_05539_),
    .ZN(_05541_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11281_ (.A1(_02903_),
    .A2(_05535_),
    .B(_05541_),
    .ZN(_01348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11282_ (.A1(\u_cpu.rf_ram.memory[89][4] ),
    .A2(_05539_),
    .ZN(_05542_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11283_ (.A1(_02906_),
    .A2(_05535_),
    .B(_05542_),
    .ZN(_01349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11284_ (.A1(\u_cpu.rf_ram.memory[89][5] ),
    .A2(_05539_),
    .ZN(_05543_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11285_ (.A1(_02909_),
    .A2(_05536_),
    .B(_05543_),
    .ZN(_01350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11286_ (.A1(\u_cpu.rf_ram.memory[89][6] ),
    .A2(_05539_),
    .ZN(_05544_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11287_ (.A1(_02912_),
    .A2(_05536_),
    .B(_05544_),
    .ZN(_01351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11288_ (.A1(\u_cpu.rf_ram.memory[89][7] ),
    .A2(_05534_),
    .ZN(_05545_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11289_ (.A1(_02915_),
    .A2(_05536_),
    .B(_05545_),
    .ZN(_01352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11290_ (.A1(_02789_),
    .A2(_02877_),
    .ZN(_05546_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11291_ (.I(_05546_),
    .Z(_05547_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11292_ (.I(_05546_),
    .Z(_05548_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11293_ (.A1(\u_cpu.rf_ram.memory[23][0] ),
    .A2(_05548_),
    .ZN(_05549_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11294_ (.A1(_02888_),
    .A2(_05547_),
    .B(_05549_),
    .ZN(_01353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11295_ (.A1(\u_cpu.rf_ram.memory[23][1] ),
    .A2(_05548_),
    .ZN(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11296_ (.A1(_02896_),
    .A2(_05547_),
    .B(_05550_),
    .ZN(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11297_ (.I(_05546_),
    .Z(_05551_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11298_ (.A1(\u_cpu.rf_ram.memory[23][2] ),
    .A2(_05551_),
    .ZN(_05552_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11299_ (.A1(_02899_),
    .A2(_05547_),
    .B(_05552_),
    .ZN(_01355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11300_ (.A1(\u_cpu.rf_ram.memory[23][3] ),
    .A2(_05551_),
    .ZN(_05553_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11301_ (.A1(_02903_),
    .A2(_05547_),
    .B(_05553_),
    .ZN(_01356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11302_ (.A1(\u_cpu.rf_ram.memory[23][4] ),
    .A2(_05551_),
    .ZN(_05554_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11303_ (.A1(_02906_),
    .A2(_05547_),
    .B(_05554_),
    .ZN(_01357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11304_ (.A1(\u_cpu.rf_ram.memory[23][5] ),
    .A2(_05551_),
    .ZN(_05555_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11305_ (.A1(_02909_),
    .A2(_05548_),
    .B(_05555_),
    .ZN(_01358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11306_ (.A1(\u_cpu.rf_ram.memory[23][6] ),
    .A2(_05551_),
    .ZN(_05556_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11307_ (.A1(_02912_),
    .A2(_05548_),
    .B(_05556_),
    .ZN(_01359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11308_ (.A1(\u_cpu.rf_ram.memory[23][7] ),
    .A2(_05546_),
    .ZN(_05557_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11309_ (.A1(_02915_),
    .A2(_05548_),
    .B(_05557_),
    .ZN(_01360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11310_ (.A1(_04511_),
    .A2(_04037_),
    .ZN(_05558_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11311_ (.A1(\u_cpu.cpu.state.ibus_cyc ),
    .A2(_05558_),
    .ZN(_05559_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11312_ (.A1(_04907_),
    .A2(_05558_),
    .B(_05559_),
    .ZN(_01361_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _11313_ (.A1(_02648_),
    .A2(_02650_),
    .A3(\u_cpu.rf_ram.rdata[7] ),
    .Z(_05560_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11314_ (.I(_05560_),
    .Z(_01362_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _11315_ (.A1(_02648_),
    .A2(\u_cpu.rf_ram.rdata[7] ),
    .A3(\u_cpu.rf_ram_if.rtrig0 ),
    .Z(_05561_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11316_ (.I(_05561_),
    .Z(_01363_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11317_ (.A1(_04032_),
    .A2(\u_cpu.rf_ram_if.rreq_r ),
    .Z(_05562_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11318_ (.I(_05562_),
    .Z(_01364_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11319_ (.A1(\u_cpu.rf_ram_if.rcnt[1] ),
    .A2(_02717_),
    .Z(_05563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11320_ (.A1(_03119_),
    .A2(_05563_),
    .ZN(_05564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11321_ (.A1(_03134_),
    .A2(_05564_),
    .ZN(_01365_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11322_ (.D(_00026_),
    .CLK(net185),
    .Q(\u_cpu.rf_ram.memory[82][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11323_ (.D(_00027_),
    .CLK(net185),
    .Q(\u_cpu.rf_ram.memory[82][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11324_ (.D(_00028_),
    .CLK(net174),
    .Q(\u_cpu.rf_ram.memory[82][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11325_ (.D(_00029_),
    .CLK(net101),
    .Q(\u_cpu.rf_ram.memory[82][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11326_ (.D(_00030_),
    .CLK(net91),
    .Q(\u_cpu.rf_ram.memory[82][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11327_ (.D(_00031_),
    .CLK(net170),
    .Q(\u_cpu.rf_ram.memory[82][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11328_ (.D(_00032_),
    .CLK(net204),
    .Q(\u_cpu.rf_ram.memory[82][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11329_ (.D(_00033_),
    .CLK(net217),
    .Q(\u_cpu.rf_ram.memory[82][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11330_ (.D(_00034_),
    .CLK(net68),
    .Q(\u_cpu.rf_ram.memory[21][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11331_ (.D(_00035_),
    .CLK(net68),
    .Q(\u_cpu.rf_ram.memory[21][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11332_ (.D(_00036_),
    .CLK(net59),
    .Q(\u_cpu.rf_ram.memory[21][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11333_ (.D(_00037_),
    .CLK(net59),
    .Q(\u_cpu.rf_ram.memory[21][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11334_ (.D(_00038_),
    .CLK(net60),
    .Q(\u_cpu.rf_ram.memory[21][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11335_ (.D(_00039_),
    .CLK(net98),
    .Q(\u_cpu.rf_ram.memory[21][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11336_ (.D(_00040_),
    .CLK(net98),
    .Q(\u_cpu.rf_ram.memory[21][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11337_ (.D(_00041_),
    .CLK(net95),
    .Q(\u_cpu.rf_ram.memory[21][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11338_ (.D(_00042_),
    .CLK(net187),
    .Q(\u_cpu.rf_ram.memory[81][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11339_ (.D(_00043_),
    .CLK(net187),
    .Q(\u_cpu.rf_ram.memory[81][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11340_ (.D(_00044_),
    .CLK(net174),
    .Q(\u_cpu.rf_ram.memory[81][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11341_ (.D(_00045_),
    .CLK(net174),
    .Q(\u_cpu.rf_ram.memory[81][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11342_ (.D(_00046_),
    .CLK(net174),
    .Q(\u_cpu.rf_ram.memory[81][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11343_ (.D(_00047_),
    .CLK(net170),
    .Q(\u_cpu.rf_ram.memory[81][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11344_ (.D(_00048_),
    .CLK(net207),
    .Q(\u_cpu.rf_ram.memory[81][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11345_ (.D(_00049_),
    .CLK(net217),
    .Q(\u_cpu.rf_ram.memory[81][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11346_ (.D(_00050_),
    .CLK(net98),
    .Q(\u_cpu.rf_ram.memory[18][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11347_ (.D(_00051_),
    .CLK(net69),
    .Q(\u_cpu.rf_ram.memory[18][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11348_ (.D(_00052_),
    .CLK(net67),
    .Q(\u_cpu.rf_ram.memory[18][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11349_ (.D(_00053_),
    .CLK(net69),
    .Q(\u_cpu.rf_ram.memory[18][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11350_ (.D(_00054_),
    .CLK(net67),
    .Q(\u_cpu.rf_ram.memory[18][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11351_ (.D(_00055_),
    .CLK(net69),
    .Q(\u_cpu.rf_ram.memory[18][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11352_ (.D(_00056_),
    .CLK(net69),
    .Q(\u_cpu.rf_ram.memory[18][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11353_ (.D(_00057_),
    .CLK(net98),
    .Q(\u_cpu.rf_ram.memory[18][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11354_ (.D(_00058_),
    .CLK(net67),
    .Q(\u_cpu.rf_ram.memory[20][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11355_ (.D(_00059_),
    .CLK(net68),
    .Q(\u_cpu.rf_ram.memory[20][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11356_ (.D(_00060_),
    .CLK(net56),
    .Q(\u_cpu.rf_ram.memory[20][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11357_ (.D(_00061_),
    .CLK(net56),
    .Q(\u_cpu.rf_ram.memory[20][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11358_ (.D(_00062_),
    .CLK(net59),
    .Q(\u_cpu.rf_ram.memory[20][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11359_ (.D(_00063_),
    .CLK(net68),
    .Q(\u_cpu.rf_ram.memory[20][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11360_ (.D(_00064_),
    .CLK(net68),
    .Q(\u_cpu.rf_ram.memory[20][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11361_ (.D(_00065_),
    .CLK(net65),
    .Q(\u_cpu.rf_ram.memory[20][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11362_ (.D(_00066_),
    .CLK(net112),
    .Q(\u_cpu.rf_ram.memory[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11363_ (.D(_00067_),
    .CLK(net114),
    .Q(\u_cpu.rf_ram.memory[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11364_ (.D(_00068_),
    .CLK(net112),
    .Q(\u_cpu.rf_ram.memory[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11365_ (.D(_00069_),
    .CLK(net121),
    .Q(\u_cpu.rf_ram.memory[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11366_ (.D(_00070_),
    .CLK(net122),
    .Q(\u_cpu.rf_ram.memory[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11367_ (.D(_00071_),
    .CLK(net123),
    .Q(\u_cpu.rf_ram.memory[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11368_ (.D(_00072_),
    .CLK(net134),
    .Q(\u_cpu.rf_ram.memory[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11369_ (.D(_00073_),
    .CLK(net133),
    .Q(\u_cpu.rf_ram.memory[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11370_ (.D(_00074_),
    .CLK(net110),
    .Q(\u_cpu.rf_ram.memory[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11371_ (.D(_00075_),
    .CLK(net114),
    .Q(\u_cpu.rf_ram.memory[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11372_ (.D(_00076_),
    .CLK(net110),
    .Q(\u_cpu.rf_ram.memory[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11373_ (.D(_00077_),
    .CLK(net60),
    .Q(\u_cpu.rf_ram.memory[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11374_ (.D(_00078_),
    .CLK(net121),
    .Q(\u_cpu.rf_ram.memory[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11375_ (.D(_00079_),
    .CLK(net122),
    .Q(\u_cpu.rf_ram.memory[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11376_ (.D(_00080_),
    .CLK(net134),
    .Q(\u_cpu.rf_ram.memory[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11377_ (.D(_00081_),
    .CLK(net133),
    .Q(\u_cpu.rf_ram.memory[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11378_ (.D(_00082_),
    .CLK(net187),
    .Q(\u_cpu.rf_ram.memory[80][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11379_ (.D(_00083_),
    .CLK(net215),
    .Q(\u_cpu.rf_ram.memory[80][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11380_ (.D(_00084_),
    .CLK(net176),
    .Q(\u_cpu.rf_ram.memory[80][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11381_ (.D(_00085_),
    .CLK(net176),
    .Q(\u_cpu.rf_ram.memory[80][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11382_ (.D(_00086_),
    .CLK(net185),
    .Q(\u_cpu.rf_ram.memory[80][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11383_ (.D(_00087_),
    .CLK(net215),
    .Q(\u_cpu.rf_ram.memory[80][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11384_ (.D(_00088_),
    .CLK(net217),
    .Q(\u_cpu.rf_ram.memory[80][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11385_ (.D(_00089_),
    .CLK(net217),
    .Q(\u_cpu.rf_ram.memory[80][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11386_ (.D(_00090_),
    .CLK(net220),
    .Q(\u_cpu.rf_ram.memory[78][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11387_ (.D(_00091_),
    .CLK(net220),
    .Q(\u_cpu.rf_ram.memory[78][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11388_ (.D(_00092_),
    .CLK(net188),
    .Q(\u_cpu.rf_ram.memory[78][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11389_ (.D(_00093_),
    .CLK(net182),
    .Q(\u_cpu.rf_ram.memory[78][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11390_ (.D(_00094_),
    .CLK(net189),
    .Q(\u_cpu.rf_ram.memory[78][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11391_ (.D(_00095_),
    .CLK(net190),
    .Q(\u_cpu.rf_ram.memory[78][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11392_ (.D(_00096_),
    .CLK(net221),
    .Q(\u_cpu.rf_ram.memory[78][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11393_ (.D(_00097_),
    .CLK(net249),
    .Q(\u_cpu.rf_ram.memory[78][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11394_ (.D(_00098_),
    .CLK(net297),
    .Q(\u_cpu.rf_ram.memory[42][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11395_ (.D(_00099_),
    .CLK(net295),
    .Q(\u_cpu.rf_ram.memory[42][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11396_ (.D(_00100_),
    .CLK(net302),
    .Q(\u_cpu.rf_ram.memory[42][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11397_ (.D(_00101_),
    .CLK(net299),
    .Q(\u_cpu.rf_ram.memory[42][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11398_ (.D(_00102_),
    .CLK(net301),
    .Q(\u_cpu.rf_ram.memory[42][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11399_ (.D(_00103_),
    .CLK(net293),
    .Q(\u_cpu.rf_ram.memory[42][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11400_ (.D(_00104_),
    .CLK(net293),
    .Q(\u_cpu.rf_ram.memory[42][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11401_ (.D(_00105_),
    .CLK(net294),
    .Q(\u_cpu.rf_ram.memory[42][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11402_ (.D(_00106_),
    .CLK(net217),
    .Q(\u_cpu.rf_ram.memory[46][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11403_ (.D(_00107_),
    .CLK(net218),
    .Q(\u_cpu.rf_ram.memory[46][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11404_ (.D(_00108_),
    .CLK(net221),
    .Q(\u_cpu.rf_ram.memory[46][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11405_ (.D(_00109_),
    .CLK(net221),
    .Q(\u_cpu.rf_ram.memory[46][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11406_ (.D(_00110_),
    .CLK(net221),
    .Q(\u_cpu.rf_ram.memory[46][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11407_ (.D(_00111_),
    .CLK(net218),
    .Q(\u_cpu.rf_ram.memory[46][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11408_ (.D(_00112_),
    .CLK(net224),
    .Q(\u_cpu.rf_ram.memory[46][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11409_ (.D(_00113_),
    .CLK(net224),
    .Q(\u_cpu.rf_ram.memory[46][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11410_ (.D(_00114_),
    .CLK(net224),
    .Q(\u_cpu.rf_ram.memory[45][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11411_ (.D(_00115_),
    .CLK(net224),
    .Q(\u_cpu.rf_ram.memory[45][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11412_ (.D(_00116_),
    .CLK(net226),
    .Q(\u_cpu.rf_ram.memory[45][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11413_ (.D(_00117_),
    .CLK(net227),
    .Q(\u_cpu.rf_ram.memory[45][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11414_ (.D(_00118_),
    .CLK(net226),
    .Q(\u_cpu.rf_ram.memory[45][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11415_ (.D(_00119_),
    .CLK(net224),
    .Q(\u_cpu.rf_ram.memory[45][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11416_ (.D(_00120_),
    .CLK(net225),
    .Q(\u_cpu.rf_ram.memory[45][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11417_ (.D(_00121_),
    .CLK(net225),
    .Q(\u_cpu.rf_ram.memory[45][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11418_ (.D(_00122_),
    .CLK(net291),
    .Q(\u_cpu.rf_ram.memory[44][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11419_ (.D(_00123_),
    .CLK(net291),
    .Q(\u_cpu.rf_ram.memory[44][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11420_ (.D(_00124_),
    .CLK(net297),
    .Q(\u_cpu.rf_ram.memory[44][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11421_ (.D(_00125_),
    .CLK(net297),
    .Q(\u_cpu.rf_ram.memory[44][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11422_ (.D(_00126_),
    .CLK(net291),
    .Q(\u_cpu.rf_ram.memory[44][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11423_ (.D(_00127_),
    .CLK(net292),
    .Q(\u_cpu.rf_ram.memory[44][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11424_ (.D(_00128_),
    .CLK(net292),
    .Q(\u_cpu.rf_ram.memory[44][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11425_ (.D(_00129_),
    .CLK(net291),
    .Q(\u_cpu.rf_ram.memory[44][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11426_ (.D(_00130_),
    .CLK(net326),
    .Q(\u_cpu.rf_ram.memory[51][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11427_ (.D(_00131_),
    .CLK(net420),
    .Q(\u_cpu.rf_ram.memory[51][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11428_ (.D(_00132_),
    .CLK(net333),
    .Q(\u_cpu.rf_ram.memory[51][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11429_ (.D(_00133_),
    .CLK(net327),
    .Q(\u_cpu.rf_ram.memory[51][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11430_ (.D(_00134_),
    .CLK(net370),
    .Q(\u_cpu.rf_ram.memory[51][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11431_ (.D(_00135_),
    .CLK(net368),
    .Q(\u_cpu.rf_ram.memory[51][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11432_ (.D(_00136_),
    .CLK(net368),
    .Q(\u_cpu.rf_ram.memory[51][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11433_ (.D(_00137_),
    .CLK(net326),
    .Q(\u_cpu.rf_ram.memory[51][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11434_ (.D(_00138_),
    .CLK(net327),
    .Q(\u_cpu.rf_ram.memory[41][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11435_ (.D(_00139_),
    .CLK(net334),
    .Q(\u_cpu.rf_ram.memory[41][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11436_ (.D(_00140_),
    .CLK(net327),
    .Q(\u_cpu.rf_ram.memory[41][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11437_ (.D(_00141_),
    .CLK(net324),
    .Q(\u_cpu.rf_ram.memory[41][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11438_ (.D(_00142_),
    .CLK(net330),
    .Q(\u_cpu.rf_ram.memory[41][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11439_ (.D(_00143_),
    .CLK(net330),
    .Q(\u_cpu.rf_ram.memory[41][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11440_ (.D(_00144_),
    .CLK(net324),
    .Q(\u_cpu.rf_ram.memory[41][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11441_ (.D(_00145_),
    .CLK(net325),
    .Q(\u_cpu.rf_ram.memory[41][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11442_ (.D(_00146_),
    .CLK(net295),
    .Q(\u_cpu.rf_ram.memory[43][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11443_ (.D(_00147_),
    .CLK(net295),
    .Q(\u_cpu.rf_ram.memory[43][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11444_ (.D(_00148_),
    .CLK(net326),
    .Q(\u_cpu.rf_ram.memory[43][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11445_ (.D(_00149_),
    .CLK(net325),
    .Q(\u_cpu.rf_ram.memory[43][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11446_ (.D(_00150_),
    .CLK(net326),
    .Q(\u_cpu.rf_ram.memory[43][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11447_ (.D(_00151_),
    .CLK(net300),
    .Q(\u_cpu.rf_ram.memory[43][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11448_ (.D(_00152_),
    .CLK(net299),
    .Q(\u_cpu.rf_ram.memory[43][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11449_ (.D(_00153_),
    .CLK(net299),
    .Q(\u_cpu.rf_ram.memory[43][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11450_ (.D(_00154_),
    .CLK(net334),
    .Q(\u_cpu.rf_ram.memory[48][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11451_ (.D(_00155_),
    .CLK(net333),
    .Q(\u_cpu.rf_ram.memory[48][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11452_ (.D(_00156_),
    .CLK(net335),
    .Q(\u_cpu.rf_ram.memory[48][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11453_ (.D(_00157_),
    .CLK(net334),
    .Q(\u_cpu.rf_ram.memory[48][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11454_ (.D(_00158_),
    .CLK(net334),
    .Q(\u_cpu.rf_ram.memory[48][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11455_ (.D(_00159_),
    .CLK(net370),
    .Q(\u_cpu.rf_ram.memory[48][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11456_ (.D(_00160_),
    .CLK(net370),
    .Q(\u_cpu.rf_ram.memory[48][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11457_ (.D(_00161_),
    .CLK(net327),
    .Q(\u_cpu.rf_ram.memory[48][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11458_ (.D(_00162_),
    .CLK(net222),
    .Q(\u_cpu.rf_ram.memory[47][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11459_ (.D(_00163_),
    .CLK(net222),
    .Q(\u_cpu.rf_ram.memory[47][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11460_ (.D(_00164_),
    .CLK(net227),
    .Q(\u_cpu.rf_ram.memory[47][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11461_ (.D(_00165_),
    .CLK(net227),
    .Q(\u_cpu.rf_ram.memory[47][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11462_ (.D(_00166_),
    .CLK(net297),
    .Q(\u_cpu.rf_ram.memory[47][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11463_ (.D(_00167_),
    .CLK(net226),
    .Q(\u_cpu.rf_ram.memory[47][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11464_ (.D(_00168_),
    .CLK(net226),
    .Q(\u_cpu.rf_ram.memory[47][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11465_ (.D(_00169_),
    .CLK(net226),
    .Q(\u_cpu.rf_ram.memory[47][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11466_ (.D(_00170_),
    .CLK(net301),
    .Q(\u_cpu.rf_ram.memory[50][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11467_ (.D(_00171_),
    .CLK(net301),
    .Q(\u_cpu.rf_ram.memory[50][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11468_ (.D(_00172_),
    .CLK(net302),
    .Q(\u_cpu.rf_ram.memory[50][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11469_ (.D(_00173_),
    .CLK(net302),
    .Q(\u_cpu.rf_ram.memory[50][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11470_ (.D(_00174_),
    .CLK(net347),
    .Q(\u_cpu.rf_ram.memory[50][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11471_ (.D(_00175_),
    .CLK(net346),
    .Q(\u_cpu.rf_ram.memory[50][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11472_ (.D(_00176_),
    .CLK(net346),
    .Q(\u_cpu.rf_ram.memory[50][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11473_ (.D(_00177_),
    .CLK(net303),
    .Q(\u_cpu.rf_ram.memory[50][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11474_ (.D(_00178_),
    .CLK(net110),
    .Q(\u_cpu.rf_ram.memory[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11475_ (.D(_00179_),
    .CLK(net121),
    .Q(\u_cpu.rf_ram.memory[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11476_ (.D(_00180_),
    .CLK(net111),
    .Q(\u_cpu.rf_ram.memory[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11477_ (.D(_00181_),
    .CLK(net67),
    .Q(\u_cpu.rf_ram.memory[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11478_ (.D(_00182_),
    .CLK(net121),
    .Q(\u_cpu.rf_ram.memory[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11479_ (.D(_00183_),
    .CLK(net122),
    .Q(\u_cpu.rf_ram.memory[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11480_ (.D(_00184_),
    .CLK(net142),
    .Q(\u_cpu.rf_ram.memory[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11481_ (.D(_00185_),
    .CLK(net133),
    .Q(\u_cpu.rf_ram.memory[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11482_ (.D(_00186_),
    .CLK(net379),
    .Q(\u_cpu.rf_ram_if.rreq_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11483_ (.D(_00187_),
    .CLK(net378),
    .Q(\u_cpu.rf_ram_if.rcnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11484_ (.D(_00188_),
    .CLK(net378),
    .Q(\u_cpu.rf_ram_if.rcnt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11485_ (.D(_00189_),
    .CLK(net376),
    .Q(\u_cpu.raddr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11486_ (.D(_00190_),
    .CLK(net376),
    .Q(\u_cpu.raddr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11487_ (.D(_00191_),
    .CLK(net99),
    .Q(\u_cpu.rf_ram.memory[16][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11488_ (.D(_00192_),
    .CLK(net105),
    .Q(\u_cpu.rf_ram.memory[16][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11489_ (.D(_00193_),
    .CLK(net178),
    .Q(\u_cpu.rf_ram.memory[16][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11490_ (.D(_00194_),
    .CLK(net178),
    .Q(\u_cpu.rf_ram.memory[16][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11491_ (.D(_00195_),
    .CLK(net180),
    .Q(\u_cpu.rf_ram.memory[16][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11492_ (.D(_00196_),
    .CLK(net105),
    .Q(\u_cpu.rf_ram.memory[16][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11493_ (.D(_00197_),
    .CLK(net105),
    .Q(\u_cpu.rf_ram.memory[16][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11494_ (.D(_00198_),
    .CLK(net98),
    .Q(\u_cpu.rf_ram.memory[16][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11495_ (.D(_00199_),
    .CLK(net99),
    .Q(\u_cpu.rf_ram.memory[17][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11496_ (.D(_00200_),
    .CLK(net140),
    .Q(\u_cpu.rf_ram.memory[17][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11497_ (.D(_00201_),
    .CLK(net178),
    .Q(\u_cpu.rf_ram.memory[17][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11498_ (.D(_00202_),
    .CLK(net178),
    .Q(\u_cpu.rf_ram.memory[17][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11499_ (.D(_00203_),
    .CLK(net178),
    .Q(\u_cpu.rf_ram.memory[17][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11500_ (.D(_00204_),
    .CLK(net106),
    .Q(\u_cpu.rf_ram.memory[17][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11501_ (.D(_00205_),
    .CLK(net106),
    .Q(\u_cpu.rf_ram.memory[17][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11502_ (.D(_00206_),
    .CLK(net99),
    .Q(\u_cpu.rf_ram.memory[17][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11503_ (.D(_00207_),
    .CLK(net295),
    .Q(\u_cpu.rf_ram.memory[40][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11504_ (.D(_00208_),
    .CLK(net295),
    .Q(\u_cpu.rf_ram.memory[40][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11505_ (.D(_00209_),
    .CLK(net302),
    .Q(\u_cpu.rf_ram.memory[40][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11506_ (.D(_00210_),
    .CLK(net326),
    .Q(\u_cpu.rf_ram.memory[40][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11507_ (.D(_00211_),
    .CLK(net302),
    .Q(\u_cpu.rf_ram.memory[40][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11508_ (.D(_00212_),
    .CLK(net303),
    .Q(\u_cpu.rf_ram.memory[40][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11509_ (.D(_00213_),
    .CLK(net301),
    .Q(\u_cpu.rf_ram.memory[40][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11510_ (.D(_00214_),
    .CLK(net301),
    .Q(\u_cpu.rf_ram.memory[40][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11511_ (.D(_00215_),
    .CLK(net320),
    .Q(\u_cpu.rf_ram.memory[119][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11512_ (.D(_00216_),
    .CLK(net319),
    .Q(\u_cpu.rf_ram.memory[119][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11513_ (.D(_00217_),
    .CLK(net320),
    .Q(\u_cpu.rf_ram.memory[119][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11514_ (.D(_00218_),
    .CLK(net320),
    .Q(\u_cpu.rf_ram.memory[119][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11515_ (.D(_00219_),
    .CLK(net321),
    .Q(\u_cpu.rf_ram.memory[119][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11516_ (.D(_00220_),
    .CLK(net400),
    .Q(\u_cpu.rf_ram.memory[119][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11517_ (.D(_00221_),
    .CLK(net400),
    .Q(\u_cpu.rf_ram.memory[119][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11518_ (.D(_00222_),
    .CLK(net321),
    .Q(\u_cpu.rf_ram.memory[119][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11519_ (.D(_00223_),
    .CLK(net430),
    .Q(\u_cpu.rf_ram.memory[129][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11520_ (.D(_00224_),
    .CLK(net430),
    .Q(\u_cpu.rf_ram.memory[129][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11521_ (.D(_00225_),
    .CLK(net430),
    .Q(\u_cpu.rf_ram.memory[129][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11522_ (.D(_00226_),
    .CLK(net430),
    .Q(\u_cpu.rf_ram.memory[129][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11523_ (.D(_00227_),
    .CLK(net431),
    .Q(\u_cpu.rf_ram.memory[129][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11524_ (.D(_00228_),
    .CLK(net432),
    .Q(\u_cpu.rf_ram.memory[129][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11525_ (.D(_00229_),
    .CLK(net430),
    .Q(\u_cpu.rf_ram.memory[129][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11526_ (.D(_00230_),
    .CLK(net432),
    .Q(\u_cpu.rf_ram.memory[129][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11527_ (.D(_00231_),
    .CLK(net488),
    .Q(\u_cpu.rf_ram.memory[139][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11528_ (.D(_00232_),
    .CLK(net511),
    .Q(\u_cpu.rf_ram.memory[139][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11529_ (.D(_00233_),
    .CLK(net488),
    .Q(\u_cpu.rf_ram.memory[139][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11530_ (.D(_00234_),
    .CLK(net488),
    .Q(\u_cpu.rf_ram.memory[139][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11531_ (.D(_00235_),
    .CLK(net489),
    .Q(\u_cpu.rf_ram.memory[139][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11532_ (.D(_00236_),
    .CLK(net486),
    .Q(\u_cpu.rf_ram.memory[139][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11533_ (.D(_00237_),
    .CLK(net488),
    .Q(\u_cpu.rf_ram.memory[139][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11534_ (.D(_00238_),
    .CLK(net488),
    .Q(\u_cpu.rf_ram.memory[139][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11535_ (.D(_00239_),
    .CLK(net250),
    .Q(\u_cpu.rf_ram.memory[77][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11536_ (.D(_00240_),
    .CLK(net250),
    .Q(\u_cpu.rf_ram.memory[77][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11537_ (.D(_00241_),
    .CLK(net241),
    .Q(\u_cpu.rf_ram.memory[77][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11538_ (.D(_00242_),
    .CLK(net234),
    .Q(\u_cpu.rf_ram.memory[77][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11539_ (.D(_00243_),
    .CLK(net242),
    .Q(\u_cpu.rf_ram.memory[77][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11540_ (.D(_00244_),
    .CLK(net249),
    .Q(\u_cpu.rf_ram.memory[77][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11541_ (.D(_00245_),
    .CLK(net249),
    .Q(\u_cpu.rf_ram.memory[77][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11542_ (.D(_00246_),
    .CLK(net250),
    .Q(\u_cpu.rf_ram.memory[77][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11543_ (.D(_00247_),
    .CLK(net256),
    .Q(\u_cpu.rf_ram.memory[74][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11544_ (.D(_00248_),
    .CLK(net261),
    .Q(\u_cpu.rf_ram.memory[74][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11545_ (.D(_00249_),
    .CLK(net258),
    .Q(\u_cpu.rf_ram.memory[74][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11546_ (.D(_00250_),
    .CLK(net258),
    .Q(\u_cpu.rf_ram.memory[74][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11547_ (.D(_00251_),
    .CLK(net258),
    .Q(\u_cpu.rf_ram.memory[74][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11548_ (.D(_00252_),
    .CLK(net339),
    .Q(\u_cpu.rf_ram.memory[74][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11549_ (.D(_00253_),
    .CLK(net339),
    .Q(\u_cpu.rf_ram.memory[74][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11550_ (.D(_00254_),
    .CLK(net261),
    .Q(\u_cpu.rf_ram.memory[74][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11551_ (.D(_00255_),
    .CLK(net250),
    .Q(\u_cpu.rf_ram.memory[76][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11552_ (.D(_00256_),
    .CLK(net253),
    .Q(\u_cpu.rf_ram.memory[76][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11553_ (.D(_00257_),
    .CLK(net241),
    .Q(\u_cpu.rf_ram.memory[76][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11554_ (.D(_00258_),
    .CLK(net241),
    .Q(\u_cpu.rf_ram.memory[76][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11555_ (.D(_00259_),
    .CLK(net242),
    .Q(\u_cpu.rf_ram.memory[76][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11556_ (.D(_00260_),
    .CLK(net249),
    .Q(\u_cpu.rf_ram.memory[76][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11557_ (.D(_00261_),
    .CLK(net249),
    .Q(\u_cpu.rf_ram.memory[76][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11558_ (.D(_00262_),
    .CLK(net250),
    .Q(\u_cpu.rf_ram.memory[76][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11559_ (.D(_00263_),
    .CLK(net257),
    .Q(\u_cpu.rf_ram.memory[75][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11560_ (.D(_00264_),
    .CLK(net258),
    .Q(\u_cpu.rf_ram.memory[75][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11561_ (.D(_00265_),
    .CLK(net258),
    .Q(\u_cpu.rf_ram.memory[75][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11562_ (.D(_00266_),
    .CLK(net259),
    .Q(\u_cpu.rf_ram.memory[75][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11563_ (.D(_00267_),
    .CLK(net341),
    .Q(\u_cpu.rf_ram.memory[75][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11564_ (.D(_00268_),
    .CLK(net343),
    .Q(\u_cpu.rf_ram.memory[75][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11565_ (.D(_00269_),
    .CLK(net341),
    .Q(\u_cpu.rf_ram.memory[75][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11566_ (.D(_00270_),
    .CLK(net341),
    .Q(\u_cpu.rf_ram.memory[75][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11567_ (.D(_00271_),
    .CLK(net110),
    .Q(\u_cpu.rf_ram.memory[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11568_ (.D(_00272_),
    .CLK(net114),
    .Q(\u_cpu.rf_ram.memory[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11569_ (.D(_00273_),
    .CLK(net110),
    .Q(\u_cpu.rf_ram.memory[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11570_ (.D(_00274_),
    .CLK(net60),
    .Q(\u_cpu.rf_ram.memory[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11571_ (.D(_00275_),
    .CLK(net114),
    .Q(\u_cpu.rf_ram.memory[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11572_ (.D(_00276_),
    .CLK(net122),
    .Q(\u_cpu.rf_ram.memory[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11573_ (.D(_00277_),
    .CLK(net134),
    .Q(\u_cpu.rf_ram.memory[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11574_ (.D(_00278_),
    .CLK(net133),
    .Q(\u_cpu.rf_ram.memory[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11575_ (.D(_00279_),
    .CLK(net340),
    .Q(\u_cpu.rf_ram.memory[68][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11576_ (.D(_00280_),
    .CLK(net340),
    .Q(\u_cpu.rf_ram.memory[68][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11577_ (.D(_00281_),
    .CLK(net347),
    .Q(\u_cpu.rf_ram.memory[68][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11578_ (.D(_00282_),
    .CLK(net349),
    .Q(\u_cpu.rf_ram.memory[68][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11579_ (.D(_00283_),
    .CLK(net350),
    .Q(\u_cpu.rf_ram.memory[68][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11580_ (.D(_00284_),
    .CLK(net340),
    .Q(\u_cpu.rf_ram.memory[68][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11581_ (.D(_00285_),
    .CLK(net339),
    .Q(\u_cpu.rf_ram.memory[68][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11582_ (.D(_00286_),
    .CLK(net340),
    .Q(\u_cpu.rf_ram.memory[68][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11583_ (.D(_00287_),
    .CLK(net245),
    .Q(\u_cpu.rf_ram.memory[67][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11584_ (.D(_00288_),
    .CLK(net245),
    .Q(\u_cpu.rf_ram.memory[67][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11585_ (.D(_00289_),
    .CLK(net248),
    .Q(\u_cpu.rf_ram.memory[67][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11586_ (.D(_00290_),
    .CLK(net248),
    .Q(\u_cpu.rf_ram.memory[67][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11587_ (.D(_00291_),
    .CLK(net251),
    .Q(\u_cpu.rf_ram.memory[67][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11588_ (.D(_00292_),
    .CLK(net252),
    .Q(\u_cpu.rf_ram.memory[67][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11589_ (.D(_00293_),
    .CLK(net253),
    .Q(\u_cpu.rf_ram.memory[67][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11590_ (.D(_00294_),
    .CLK(net253),
    .Q(\u_cpu.rf_ram.memory[67][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11591_ (.D(_00295_),
    .CLK(net245),
    .Q(\u_cpu.rf_ram.memory[66][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11592_ (.D(_00296_),
    .CLK(net245),
    .Q(\u_cpu.rf_ram.memory[66][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11593_ (.D(_00297_),
    .CLK(net244),
    .Q(\u_cpu.rf_ram.memory[66][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11594_ (.D(_00298_),
    .CLK(net246),
    .Q(\u_cpu.rf_ram.memory[66][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11595_ (.D(_00299_),
    .CLK(net251),
    .Q(\u_cpu.rf_ram.memory[66][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11596_ (.D(_00300_),
    .CLK(net251),
    .Q(\u_cpu.rf_ram.memory[66][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11597_ (.D(_00301_),
    .CLK(net251),
    .Q(\u_cpu.rf_ram.memory[66][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11598_ (.D(_00302_),
    .CLK(net251),
    .Q(\u_cpu.rf_ram.memory[66][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11599_ (.D(_00303_),
    .CLK(net244),
    .Q(\u_cpu.rf_ram.memory[65][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11600_ (.D(_00304_),
    .CLK(net244),
    .Q(\u_cpu.rf_ram.memory[65][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11601_ (.D(_00305_),
    .CLK(net243),
    .Q(\u_cpu.rf_ram.memory[65][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11602_ (.D(_00306_),
    .CLK(net243),
    .Q(\u_cpu.rf_ram.memory[65][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11603_ (.D(_00307_),
    .CLK(net243),
    .Q(\u_cpu.rf_ram.memory[65][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11604_ (.D(_00308_),
    .CLK(net243),
    .Q(\u_cpu.rf_ram.memory[65][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11605_ (.D(_00309_),
    .CLK(net243),
    .Q(\u_cpu.rf_ram.memory[65][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11606_ (.D(_00310_),
    .CLK(net244),
    .Q(\u_cpu.rf_ram.memory[65][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11607_ (.D(_00311_),
    .CLK(net236),
    .Q(\u_cpu.rf_ram.memory[64][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11608_ (.D(_00312_),
    .CLK(net236),
    .Q(\u_cpu.rf_ram.memory[64][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11609_ (.D(_00313_),
    .CLK(net236),
    .Q(\u_cpu.rf_ram.memory[64][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11610_ (.D(_00314_),
    .CLK(net237),
    .Q(\u_cpu.rf_ram.memory[64][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11611_ (.D(_00315_),
    .CLK(net238),
    .Q(\u_cpu.rf_ram.memory[64][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11612_ (.D(_00316_),
    .CLK(net238),
    .Q(\u_cpu.rf_ram.memory[64][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11613_ (.D(_00317_),
    .CLK(net238),
    .Q(\u_cpu.rf_ram.memory[64][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11614_ (.D(_00318_),
    .CLK(net239),
    .Q(\u_cpu.rf_ram.memory[64][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11615_ (.D(_00319_),
    .CLK(net101),
    .Q(\u_cpu.rf_ram.memory[29][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11616_ (.D(_00320_),
    .CLK(net101),
    .Q(\u_cpu.rf_ram.memory[29][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11617_ (.D(_00321_),
    .CLK(net103),
    .Q(\u_cpu.rf_ram.memory[29][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11618_ (.D(_00322_),
    .CLK(net103),
    .Q(\u_cpu.rf_ram.memory[29][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11619_ (.D(_00323_),
    .CLK(net103),
    .Q(\u_cpu.rf_ram.memory[29][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11620_ (.D(_00324_),
    .CLK(net101),
    .Q(\u_cpu.rf_ram.memory[29][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11621_ (.D(_00325_),
    .CLK(net101),
    .Q(\u_cpu.rf_ram.memory[29][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11622_ (.D(_00326_),
    .CLK(net174),
    .Q(\u_cpu.rf_ram.memory[29][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11623_ (.D(_00327_),
    .CLK(net185),
    .Q(\u_cpu.rf_ram.memory[63][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11624_ (.D(_00328_),
    .CLK(net186),
    .Q(\u_cpu.rf_ram.memory[63][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11625_ (.D(_00329_),
    .CLK(net176),
    .Q(\u_cpu.rf_ram.memory[63][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11626_ (.D(_00330_),
    .CLK(net177),
    .Q(\u_cpu.rf_ram.memory[63][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11627_ (.D(_00331_),
    .CLK(net177),
    .Q(\u_cpu.rf_ram.memory[63][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11628_ (.D(_00332_),
    .CLK(net181),
    .Q(\u_cpu.rf_ram.memory[63][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11629_ (.D(_00333_),
    .CLK(net181),
    .Q(\u_cpu.rf_ram.memory[63][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11630_ (.D(_00334_),
    .CLK(net181),
    .Q(\u_cpu.rf_ram.memory[63][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11631_ (.D(_00335_),
    .CLK(net175),
    .Q(\u_cpu.rf_ram.memory[62][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11632_ (.D(_00336_),
    .CLK(net175),
    .Q(\u_cpu.rf_ram.memory[62][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11633_ (.D(_00337_),
    .CLK(net175),
    .Q(\u_cpu.rf_ram.memory[62][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11634_ (.D(_00338_),
    .CLK(net175),
    .Q(\u_cpu.rf_ram.memory[62][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11635_ (.D(_00339_),
    .CLK(net175),
    .Q(\u_cpu.rf_ram.memory[62][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11636_ (.D(_00340_),
    .CLK(net179),
    .Q(\u_cpu.rf_ram.memory[62][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11637_ (.D(_00341_),
    .CLK(net179),
    .Q(\u_cpu.rf_ram.memory[62][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11638_ (.D(_00342_),
    .CLK(net179),
    .Q(\u_cpu.rf_ram.memory[62][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11639_ (.D(_00343_),
    .CLK(net186),
    .Q(\u_cpu.rf_ram.memory[61][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11640_ (.D(_00344_),
    .CLK(net188),
    .Q(\u_cpu.rf_ram.memory[61][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11641_ (.D(_00345_),
    .CLK(net188),
    .Q(\u_cpu.rf_ram.memory[61][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11642_ (.D(_00346_),
    .CLK(net189),
    .Q(\u_cpu.rf_ram.memory[61][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11643_ (.D(_00347_),
    .CLK(net189),
    .Q(\u_cpu.rf_ram.memory[61][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11644_ (.D(_00348_),
    .CLK(net188),
    .Q(\u_cpu.rf_ram.memory[61][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11645_ (.D(_00349_),
    .CLK(net189),
    .Q(\u_cpu.rf_ram.memory[61][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11646_ (.D(_00350_),
    .CLK(net189),
    .Q(\u_cpu.rf_ram.memory[61][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11647_ (.D(_00351_),
    .CLK(net215),
    .Q(\u_cpu.rf_ram.memory[60][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11648_ (.D(_00352_),
    .CLK(net215),
    .Q(\u_cpu.rf_ram.memory[60][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11649_ (.D(_00353_),
    .CLK(net215),
    .Q(\u_cpu.rf_ram.memory[60][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11650_ (.D(_00354_),
    .CLK(net216),
    .Q(\u_cpu.rf_ram.memory[60][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11651_ (.D(_00355_),
    .CLK(net216),
    .Q(\u_cpu.rf_ram.memory[60][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11652_ (.D(_00356_),
    .CLK(net220),
    .Q(\u_cpu.rf_ram.memory[60][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11653_ (.D(_00357_),
    .CLK(net220),
    .Q(\u_cpu.rf_ram.memory[60][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11654_ (.D(_00358_),
    .CLK(net220),
    .Q(\u_cpu.rf_ram.memory[60][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11655_ (.D(_00359_),
    .CLK(net179),
    .Q(\u_cpu.rf_ram.memory[19][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11656_ (.D(_00360_),
    .CLK(net179),
    .Q(\u_cpu.rf_ram.memory[19][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11657_ (.D(_00361_),
    .CLK(net181),
    .Q(\u_cpu.rf_ram.memory[19][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11658_ (.D(_00362_),
    .CLK(net181),
    .Q(\u_cpu.rf_ram.memory[19][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11659_ (.D(_00363_),
    .CLK(net182),
    .Q(\u_cpu.rf_ram.memory[19][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11660_ (.D(_00364_),
    .CLK(net188),
    .Q(\u_cpu.rf_ram.memory[19][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11661_ (.D(_00365_),
    .CLK(net191),
    .Q(\u_cpu.rf_ram.memory[19][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11662_ (.D(_00366_),
    .CLK(net182),
    .Q(\u_cpu.rf_ram.memory[19][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11663_ (.D(_00367_),
    .CLK(net111),
    .Q(\u_cpu.rf_ram.memory[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11664_ (.D(_00368_),
    .CLK(net121),
    .Q(\u_cpu.rf_ram.memory[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11665_ (.D(_00369_),
    .CLK(net58),
    .Q(\u_cpu.rf_ram.memory[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11666_ (.D(_00370_),
    .CLK(net70),
    .Q(\u_cpu.rf_ram.memory[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11667_ (.D(_00371_),
    .CLK(net114),
    .Q(\u_cpu.rf_ram.memory[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11668_ (.D(_00372_),
    .CLK(net122),
    .Q(\u_cpu.rf_ram.memory[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11669_ (.D(_00373_),
    .CLK(net142),
    .Q(\u_cpu.rf_ram.memory[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11670_ (.D(_00374_),
    .CLK(net99),
    .Q(\u_cpu.rf_ram.memory[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11671_ (.D(_00375_),
    .CLK(net314),
    .Q(\u_cpu.rf_ram.memory[58][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11672_ (.D(_00376_),
    .CLK(net314),
    .Q(\u_cpu.rf_ram.memory[58][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11673_ (.D(_00377_),
    .CLK(net314),
    .Q(\u_cpu.rf_ram.memory[58][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11674_ (.D(_00378_),
    .CLK(net325),
    .Q(\u_cpu.rf_ram.memory[58][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11675_ (.D(_00379_),
    .CLK(net325),
    .Q(\u_cpu.rf_ram.memory[58][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11676_ (.D(_00380_),
    .CLK(net288),
    .Q(\u_cpu.rf_ram.memory[58][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11677_ (.D(_00381_),
    .CLK(net286),
    .Q(\u_cpu.rf_ram.memory[58][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11678_ (.D(_00382_),
    .CLK(net299),
    .Q(\u_cpu.rf_ram.memory[58][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11679_ (.D(_00383_),
    .CLK(net314),
    .Q(\u_cpu.rf_ram.memory[57][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11680_ (.D(_00384_),
    .CLK(net313),
    .Q(\u_cpu.rf_ram.memory[57][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11681_ (.D(_00385_),
    .CLK(net324),
    .Q(\u_cpu.rf_ram.memory[57][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11682_ (.D(_00386_),
    .CLK(net324),
    .Q(\u_cpu.rf_ram.memory[57][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11683_ (.D(_00387_),
    .CLK(net324),
    .Q(\u_cpu.rf_ram.memory[57][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11684_ (.D(_00388_),
    .CLK(net300),
    .Q(\u_cpu.rf_ram.memory[57][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11685_ (.D(_00389_),
    .CLK(net287),
    .Q(\u_cpu.rf_ram.memory[57][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11686_ (.D(_00390_),
    .CLK(net299),
    .Q(\u_cpu.rf_ram.memory[57][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11687_ (.D(_00391_),
    .CLK(net329),
    .Q(\u_cpu.rf_ram.memory[56][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11688_ (.D(_00392_),
    .CLK(net329),
    .Q(\u_cpu.rf_ram.memory[56][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11689_ (.D(_00393_),
    .CLK(net329),
    .Q(\u_cpu.rf_ram.memory[56][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11690_ (.D(_00394_),
    .CLK(net331),
    .Q(\u_cpu.rf_ram.memory[56][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11691_ (.D(_00395_),
    .CLK(net329),
    .Q(\u_cpu.rf_ram.memory[56][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11692_ (.D(_00396_),
    .CLK(net331),
    .Q(\u_cpu.rf_ram.memory[56][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11693_ (.D(_00397_),
    .CLK(net331),
    .Q(\u_cpu.rf_ram.memory[56][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11694_ (.D(_00398_),
    .CLK(net329),
    .Q(\u_cpu.rf_ram.memory[56][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11695_ (.D(_00399_),
    .CLK(net331),
    .Q(\u_cpu.rf_ram.memory[55][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11696_ (.D(_00400_),
    .CLK(net417),
    .Q(\u_cpu.rf_ram.memory[55][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11697_ (.D(_00401_),
    .CLK(net452),
    .Q(\u_cpu.rf_ram.memory[55][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11698_ (.D(_00402_),
    .CLK(net452),
    .Q(\u_cpu.rf_ram.memory[55][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11699_ (.D(_00403_),
    .CLK(net427),
    .Q(\u_cpu.rf_ram.memory[55][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11700_ (.D(_00404_),
    .CLK(net425),
    .Q(\u_cpu.rf_ram.memory[55][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11701_ (.D(_00405_),
    .CLK(net415),
    .Q(\u_cpu.rf_ram.memory[55][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11702_ (.D(_00406_),
    .CLK(net416),
    .Q(\u_cpu.rf_ram.memory[55][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11703_ (.D(_00407_),
    .CLK(net330),
    .Q(\u_cpu.rf_ram.memory[54][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11704_ (.D(_00408_),
    .CLK(net421),
    .Q(\u_cpu.rf_ram.memory[54][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11705_ (.D(_00409_),
    .CLK(net427),
    .Q(\u_cpu.rf_ram.memory[54][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11706_ (.D(_00410_),
    .CLK(net428),
    .Q(\u_cpu.rf_ram.memory[54][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11707_ (.D(_00411_),
    .CLK(net427),
    .Q(\u_cpu.rf_ram.memory[54][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11708_ (.D(_00412_),
    .CLK(net425),
    .Q(\u_cpu.rf_ram.memory[54][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11709_ (.D(_00413_),
    .CLK(net416),
    .Q(\u_cpu.rf_ram.memory[54][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11710_ (.D(_00414_),
    .CLK(net416),
    .Q(\u_cpu.rf_ram.memory[54][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11711_ (.D(_00415_),
    .CLK(net331),
    .Q(\u_cpu.rf_ram.memory[53][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11712_ (.D(_00416_),
    .CLK(net417),
    .Q(\u_cpu.rf_ram.memory[53][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11713_ (.D(_00417_),
    .CLK(net450),
    .Q(\u_cpu.rf_ram.memory[53][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11714_ (.D(_00418_),
    .CLK(net450),
    .Q(\u_cpu.rf_ram.memory[53][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11715_ (.D(_00419_),
    .CLK(net427),
    .Q(\u_cpu.rf_ram.memory[53][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11716_ (.D(_00420_),
    .CLK(net426),
    .Q(\u_cpu.rf_ram.memory[53][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11717_ (.D(_00421_),
    .CLK(net417),
    .Q(\u_cpu.rf_ram.memory[53][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11718_ (.D(_00422_),
    .CLK(net415),
    .Q(\u_cpu.rf_ram.memory[53][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11719_ (.D(_00423_),
    .CLK(net332),
    .Q(\u_cpu.rf_ram.memory[52][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11720_ (.D(_00424_),
    .CLK(net418),
    .Q(\u_cpu.rf_ram.memory[52][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11721_ (.D(_00425_),
    .CLK(net452),
    .Q(\u_cpu.rf_ram.memory[52][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11722_ (.D(_00426_),
    .CLK(net450),
    .Q(\u_cpu.rf_ram.memory[52][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11723_ (.D(_00427_),
    .CLK(net427),
    .Q(\u_cpu.rf_ram.memory[52][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11724_ (.D(_00428_),
    .CLK(net426),
    .Q(\u_cpu.rf_ram.memory[52][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11725_ (.D(_00429_),
    .CLK(net418),
    .Q(\u_cpu.rf_ram.memory[52][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11726_ (.D(_00430_),
    .CLK(net416),
    .Q(\u_cpu.rf_ram.memory[52][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11727_ (.D(_00431_),
    .CLK(net127),
    .Q(\u_cpu.rf_ram.memory[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11728_ (.D(_00432_),
    .CLK(net136),
    .Q(\u_cpu.rf_ram.memory[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11729_ (.D(_00433_),
    .CLK(net128),
    .Q(\u_cpu.rf_ram.memory[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11730_ (.D(_00434_),
    .CLK(net136),
    .Q(\u_cpu.rf_ram.memory[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11731_ (.D(_00435_),
    .CLK(net132),
    .Q(\u_cpu.rf_ram.memory[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11732_ (.D(_00436_),
    .CLK(net135),
    .Q(\u_cpu.rf_ram.memory[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11733_ (.D(_00437_),
    .CLK(net145),
    .Q(\u_cpu.rf_ram.memory[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11734_ (.D(_00438_),
    .CLK(net143),
    .Q(\u_cpu.rf_ram.memory[9][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11735_ (.D(_00439_),
    .CLK(net136),
    .Q(\u_cpu.rf_ram.memory[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11736_ (.D(_00440_),
    .CLK(net149),
    .Q(\u_cpu.rf_ram.memory[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11737_ (.D(_00441_),
    .CLK(net149),
    .Q(\u_cpu.rf_ram.memory[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11738_ (.D(_00442_),
    .CLK(net152),
    .Q(\u_cpu.rf_ram.memory[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11739_ (.D(_00443_),
    .CLK(net152),
    .Q(\u_cpu.rf_ram.memory[15][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11740_ (.D(_00444_),
    .CLK(net143),
    .Q(\u_cpu.rf_ram.memory[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11741_ (.D(_00445_),
    .CLK(net140),
    .Q(\u_cpu.rf_ram.memory[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11742_ (.D(_00446_),
    .CLK(net145),
    .Q(\u_cpu.rf_ram.memory[15][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11743_ (.D(_00000_),
    .CLK(net256),
    .Q(\u_cpu.rf_ram.rdata[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11744_ (.D(_00001_),
    .CLK(net252),
    .Q(\u_cpu.rf_ram.rdata[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11745_ (.D(_00002_),
    .CLK(net252),
    .Q(\u_cpu.rf_ram.rdata[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11746_ (.D(_00003_),
    .CLK(net252),
    .Q(\u_cpu.rf_ram.rdata[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11747_ (.D(_00004_),
    .CLK(net253),
    .Q(\u_cpu.rf_ram.rdata[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11748_ (.D(_00005_),
    .CLK(net256),
    .Q(\u_cpu.rf_ram.rdata[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11749_ (.D(_00006_),
    .CLK(net256),
    .Q(\u_cpu.rf_ram.rdata[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11750_ (.D(_00007_),
    .CLK(net254),
    .Q(\u_cpu.rf_ram.rdata[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11751_ (.D(_00447_),
    .CLK(net479),
    .Q(\u_cpu.rf_ram.memory[142][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11752_ (.D(_00448_),
    .CLK(net479),
    .Q(\u_cpu.rf_ram.memory[142][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11753_ (.D(_00449_),
    .CLK(net481),
    .Q(\u_cpu.rf_ram.memory[142][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11754_ (.D(_00450_),
    .CLK(net490),
    .Q(\u_cpu.rf_ram.memory[142][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11755_ (.D(_00451_),
    .CLK(net491),
    .Q(\u_cpu.rf_ram.memory[142][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11756_ (.D(_00452_),
    .CLK(net512),
    .Q(\u_cpu.rf_ram.memory[142][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11757_ (.D(_00453_),
    .CLK(net512),
    .Q(\u_cpu.rf_ram.memory[142][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11758_ (.D(_00454_),
    .CLK(net512),
    .Q(\u_cpu.rf_ram.memory[142][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11759_ (.D(_00455_),
    .CLK(net479),
    .Q(\u_cpu.rf_ram.memory[141][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11760_ (.D(_00456_),
    .CLK(net479),
    .Q(\u_cpu.rf_ram.memory[141][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11761_ (.D(_00457_),
    .CLK(net481),
    .Q(\u_cpu.rf_ram.memory[141][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11762_ (.D(_00458_),
    .CLK(net490),
    .Q(\u_cpu.rf_ram.memory[141][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11763_ (.D(_00459_),
    .CLK(net491),
    .Q(\u_cpu.rf_ram.memory[141][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11764_ (.D(_00460_),
    .CLK(net508),
    .Q(\u_cpu.rf_ram.memory[141][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11765_ (.D(_00461_),
    .CLK(net514),
    .Q(\u_cpu.rf_ram.memory[141][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11766_ (.D(_00462_),
    .CLK(net512),
    .Q(\u_cpu.rf_ram.memory[141][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11767_ (.D(_00463_),
    .CLK(net479),
    .Q(\u_cpu.rf_ram.memory[140][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11768_ (.D(_00464_),
    .CLK(net481),
    .Q(\u_cpu.rf_ram.memory[140][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11769_ (.D(_00465_),
    .CLK(net481),
    .Q(\u_cpu.rf_ram.memory[140][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11770_ (.D(_00466_),
    .CLK(net490),
    .Q(\u_cpu.rf_ram.memory[140][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11771_ (.D(_00467_),
    .CLK(net491),
    .Q(\u_cpu.rf_ram.memory[140][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11772_ (.D(_00468_),
    .CLK(net514),
    .Q(\u_cpu.rf_ram.memory[140][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11773_ (.D(_00469_),
    .CLK(net514),
    .Q(\u_cpu.rf_ram.memory[140][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11774_ (.D(_00470_),
    .CLK(net512),
    .Q(\u_cpu.rf_ram.memory[140][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11775_ (.D(_00471_),
    .CLK(net137),
    .Q(\u_cpu.rf_ram.memory[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11776_ (.D(_00472_),
    .CLK(net149),
    .Q(\u_cpu.rf_ram.memory[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11777_ (.D(_00473_),
    .CLK(net150),
    .Q(\u_cpu.rf_ram.memory[13][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11778_ (.D(_00474_),
    .CLK(net152),
    .Q(\u_cpu.rf_ram.memory[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11779_ (.D(_00475_),
    .CLK(net153),
    .Q(\u_cpu.rf_ram.memory[13][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11780_ (.D(_00476_),
    .CLK(net145),
    .Q(\u_cpu.rf_ram.memory[13][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11781_ (.D(_00477_),
    .CLK(net236),
    .Q(\u_cpu.rf_ram.memory[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11782_ (.D(_00478_),
    .CLK(net237),
    .Q(\u_cpu.rf_ram.memory[13][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11783_ (.D(_00479_),
    .CLK(net352),
    .Q(\u_cpu.rf_ram.memory[72][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11784_ (.D(_00480_),
    .CLK(net352),
    .Q(\u_cpu.rf_ram.memory[72][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11785_ (.D(_00481_),
    .CLK(net350),
    .Q(\u_cpu.rf_ram.memory[72][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11786_ (.D(_00482_),
    .CLK(net350),
    .Q(\u_cpu.rf_ram.memory[72][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11787_ (.D(_00483_),
    .CLK(net350),
    .Q(\u_cpu.rf_ram.memory[72][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11788_ (.D(_00484_),
    .CLK(net374),
    .Q(\u_cpu.rf_ram.memory[72][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11789_ (.D(_00485_),
    .CLK(net371),
    .Q(\u_cpu.rf_ram.memory[72][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11790_ (.D(_00486_),
    .CLK(net347),
    .Q(\u_cpu.rf_ram.memory[72][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11791_ (.D(_00487_),
    .CLK(net373),
    .Q(\u_cpu.rf_ram.memory[73][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11792_ (.D(_00488_),
    .CLK(net373),
    .Q(\u_cpu.rf_ram.memory[73][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11793_ (.D(_00489_),
    .CLK(net352),
    .Q(\u_cpu.rf_ram.memory[73][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11794_ (.D(_00490_),
    .CLK(net352),
    .Q(\u_cpu.rf_ram.memory[73][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11795_ (.D(_00491_),
    .CLK(net373),
    .Q(\u_cpu.rf_ram.memory[73][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11796_ (.D(_00492_),
    .CLK(net374),
    .Q(\u_cpu.rf_ram.memory[73][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11797_ (.D(_00493_),
    .CLK(net371),
    .Q(\u_cpu.rf_ram.memory[73][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11798_ (.D(_00494_),
    .CLK(net368),
    .Q(\u_cpu.rf_ram.memory[73][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11799_ (.D(_00495_),
    .CLK(net368),
    .Q(\u_cpu.rf_ram.memory[71][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11800_ (.D(_00496_),
    .CLK(net348),
    .Q(\u_cpu.rf_ram.memory[71][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11801_ (.D(_00497_),
    .CLK(net368),
    .Q(\u_cpu.rf_ram.memory[71][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11802_ (.D(_00498_),
    .CLK(net369),
    .Q(\u_cpu.rf_ram.memory[71][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11803_ (.D(_00499_),
    .CLK(net369),
    .Q(\u_cpu.rf_ram.memory[71][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11804_ (.D(_00500_),
    .CLK(net348),
    .Q(\u_cpu.rf_ram.memory[71][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11805_ (.D(_00501_),
    .CLK(net347),
    .Q(\u_cpu.rf_ram.memory[71][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11806_ (.D(_00502_),
    .CLK(net347),
    .Q(\u_cpu.rf_ram.memory[71][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11807_ (.D(_00503_),
    .CLK(net370),
    .Q(\u_cpu.rf_ram.memory[70][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11808_ (.D(_00504_),
    .CLK(net376),
    .Q(\u_cpu.rf_ram.memory[70][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11809_ (.D(_00505_),
    .CLK(net371),
    .Q(\u_cpu.rf_ram.memory[70][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11810_ (.D(_00506_),
    .CLK(net371),
    .Q(\u_cpu.rf_ram.memory[70][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11811_ (.D(_00507_),
    .CLK(net376),
    .Q(\u_cpu.rf_ram.memory[70][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11812_ (.D(_00508_),
    .CLK(net376),
    .Q(\u_cpu.rf_ram.memory[70][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11813_ (.D(_00509_),
    .CLK(net377),
    .Q(\u_cpu.rf_ram.memory[70][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11814_ (.D(_00510_),
    .CLK(net370),
    .Q(\u_cpu.rf_ram.memory[70][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11815_ (.D(_00511_),
    .CLK(net477),
    .Q(\u_cpu.rf_ram.memory[143][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11816_ (.D(_00512_),
    .CLK(net477),
    .Q(\u_cpu.rf_ram.memory[143][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11817_ (.D(_00513_),
    .CLK(net478),
    .Q(\u_cpu.rf_ram.memory[143][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11818_ (.D(_00514_),
    .CLK(net485),
    .Q(\u_cpu.rf_ram.memory[143][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11819_ (.D(_00515_),
    .CLK(net485),
    .Q(\u_cpu.rf_ram.memory[143][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11820_ (.D(_00516_),
    .CLK(net485),
    .Q(\u_cpu.rf_ram.memory[143][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11821_ (.D(_00517_),
    .CLK(net486),
    .Q(\u_cpu.rf_ram.memory[143][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11822_ (.D(_00518_),
    .CLK(net477),
    .Q(\u_cpu.rf_ram.memory[143][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11823_ (.D(_00519_),
    .CLK(net136),
    .Q(\u_cpu.rf_ram.memory[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11824_ (.D(_00520_),
    .CLK(net149),
    .Q(\u_cpu.rf_ram.memory[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11825_ (.D(_00521_),
    .CLK(net149),
    .Q(\u_cpu.rf_ram.memory[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11826_ (.D(_00522_),
    .CLK(net152),
    .Q(\u_cpu.rf_ram.memory[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11827_ (.D(_00523_),
    .CLK(net152),
    .Q(\u_cpu.rf_ram.memory[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11828_ (.D(_00524_),
    .CLK(net144),
    .Q(\u_cpu.rf_ram.memory[14][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11829_ (.D(_00525_),
    .CLK(net141),
    .Q(\u_cpu.rf_ram.memory[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11830_ (.D(_00526_),
    .CLK(net146),
    .Q(\u_cpu.rf_ram.memory[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11831_ (.D(_00527_),
    .CLK(net478),
    .Q(\u_cpu.rf_ram.memory[138][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11832_ (.D(_00528_),
    .CLK(net478),
    .Q(\u_cpu.rf_ram.memory[138][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11833_ (.D(_00529_),
    .CLK(net478),
    .Q(\u_cpu.rf_ram.memory[138][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11834_ (.D(_00530_),
    .CLK(net485),
    .Q(\u_cpu.rf_ram.memory[138][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11835_ (.D(_00531_),
    .CLK(net485),
    .Q(\u_cpu.rf_ram.memory[138][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11836_ (.D(_00532_),
    .CLK(net487),
    .Q(\u_cpu.rf_ram.memory[138][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11837_ (.D(_00533_),
    .CLK(net487),
    .Q(\u_cpu.rf_ram.memory[138][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11838_ (.D(_00534_),
    .CLK(net478),
    .Q(\u_cpu.rf_ram.memory[138][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11839_ (.D(_00535_),
    .CLK(net421),
    .Q(\u_cpu.rf_ram.memory[39][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11840_ (.D(_00536_),
    .CLK(net421),
    .Q(\u_cpu.rf_ram.memory[39][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11841_ (.D(_00537_),
    .CLK(net422),
    .Q(\u_cpu.rf_ram.memory[39][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11842_ (.D(_00538_),
    .CLK(net432),
    .Q(\u_cpu.rf_ram.memory[39][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11843_ (.D(_00539_),
    .CLK(net432),
    .Q(\u_cpu.rf_ram.memory[39][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11844_ (.D(_00540_),
    .CLK(net421),
    .Q(\u_cpu.rf_ram.memory[39][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11845_ (.D(_00541_),
    .CLK(net432),
    .Q(\u_cpu.rf_ram.memory[39][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11846_ (.D(_00542_),
    .CLK(net421),
    .Q(\u_cpu.rf_ram.memory[39][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11847_ (.D(_00543_),
    .CLK(net508),
    .Q(\u_cpu.rf_ram.memory[137][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11848_ (.D(_00544_),
    .CLK(net509),
    .Q(\u_cpu.rf_ram.memory[137][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11849_ (.D(_00545_),
    .CLK(net508),
    .Q(\u_cpu.rf_ram.memory[137][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11850_ (.D(_00546_),
    .CLK(net508),
    .Q(\u_cpu.rf_ram.memory[137][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11851_ (.D(_00547_),
    .CLK(net508),
    .Q(\u_cpu.rf_ram.memory[137][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11852_ (.D(_00548_),
    .CLK(net509),
    .Q(\u_cpu.rf_ram.memory[137][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11853_ (.D(_00549_),
    .CLK(net510),
    .Q(\u_cpu.rf_ram.memory[137][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11854_ (.D(_00550_),
    .CLK(net510),
    .Q(\u_cpu.rf_ram.memory[137][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11855_ (.D(_00551_),
    .CLK(net422),
    .Q(\u_cpu.rf_ram.memory[49][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11856_ (.D(_00552_),
    .CLK(net422),
    .Q(\u_cpu.rf_ram.memory[49][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11857_ (.D(_00553_),
    .CLK(net420),
    .Q(\u_cpu.rf_ram.memory[49][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11858_ (.D(_00554_),
    .CLK(net420),
    .Q(\u_cpu.rf_ram.memory[49][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11859_ (.D(_00555_),
    .CLK(net477),
    .Q(\u_cpu.rf_ram.memory[49][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11860_ (.D(_00556_),
    .CLK(net477),
    .Q(\u_cpu.rf_ram.memory[49][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11861_ (.D(_00557_),
    .CLK(net377),
    .Q(\u_cpu.rf_ram.memory[49][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11862_ (.D(_00558_),
    .CLK(net420),
    .Q(\u_cpu.rf_ram.memory[49][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11863_ (.D(_00559_),
    .CLK(net516),
    .Q(\u_cpu.rf_ram.memory[136][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11864_ (.D(_00560_),
    .CLK(net517),
    .Q(\u_cpu.rf_ram.memory[136][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11865_ (.D(_00561_),
    .CLK(net519),
    .Q(\u_cpu.rf_ram.memory[136][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11866_ (.D(_00562_),
    .CLK(net518),
    .Q(\u_cpu.rf_ram.memory[136][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11867_ (.D(_00563_),
    .CLK(net519),
    .Q(\u_cpu.rf_ram.memory[136][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11868_ (.D(_00564_),
    .CLK(net517),
    .Q(\u_cpu.rf_ram.memory[136][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11869_ (.D(_00565_),
    .CLK(net516),
    .Q(\u_cpu.rf_ram.memory[136][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11870_ (.D(_00566_),
    .CLK(net516),
    .Q(\u_cpu.rf_ram.memory[136][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11871_ (.D(_00567_),
    .CLK(net511),
    .Q(\u_cpu.rf_ram.memory[135][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11872_ (.D(_00568_),
    .CLK(net511),
    .Q(\u_cpu.rf_ram.memory[135][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11873_ (.D(_00569_),
    .CLK(net518),
    .Q(\u_cpu.rf_ram.memory[135][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11874_ (.D(_00570_),
    .CLK(net518),
    .Q(\u_cpu.rf_ram.memory[135][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11875_ (.D(_00571_),
    .CLK(net519),
    .Q(\u_cpu.rf_ram.memory[135][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11876_ (.D(_00572_),
    .CLK(net516),
    .Q(\u_cpu.rf_ram.memory[135][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11877_ (.D(_00573_),
    .CLK(net516),
    .Q(\u_cpu.rf_ram.memory[135][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11878_ (.D(_00574_),
    .CLK(net510),
    .Q(\u_cpu.rf_ram.memory[135][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11879_ (.D(_00575_),
    .CLK(net456),
    .Q(\u_cpu.rf_ram.memory[134][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11880_ (.D(_00576_),
    .CLK(net456),
    .Q(\u_cpu.rf_ram.memory[134][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11881_ (.D(_00577_),
    .CLK(net518),
    .Q(\u_cpu.rf_ram.memory[134][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11882_ (.D(_00578_),
    .CLK(net470),
    .Q(\u_cpu.rf_ram.memory[134][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11883_ (.D(_00579_),
    .CLK(net518),
    .Q(\u_cpu.rf_ram.memory[134][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11884_ (.D(_00580_),
    .CLK(net468),
    .Q(\u_cpu.rf_ram.memory[134][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11885_ (.D(_00581_),
    .CLK(net468),
    .Q(\u_cpu.rf_ram.memory[134][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11886_ (.D(_00582_),
    .CLK(net458),
    .Q(\u_cpu.rf_ram.memory[134][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11887_ (.D(_00583_),
    .CLK(net456),
    .Q(\u_cpu.rf_ram.memory[133][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11888_ (.D(_00584_),
    .CLK(net456),
    .Q(\u_cpu.rf_ram.memory[133][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11889_ (.D(_00585_),
    .CLK(net470),
    .Q(\u_cpu.rf_ram.memory[133][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11890_ (.D(_00586_),
    .CLK(net470),
    .Q(\u_cpu.rf_ram.memory[133][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11891_ (.D(_00587_),
    .CLK(net470),
    .Q(\u_cpu.rf_ram.memory[133][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11892_ (.D(_00588_),
    .CLK(net468),
    .Q(\u_cpu.rf_ram.memory[133][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11893_ (.D(_00589_),
    .CLK(net468),
    .Q(\u_cpu.rf_ram.memory[133][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11894_ (.D(_00590_),
    .CLK(net458),
    .Q(\u_cpu.rf_ram.memory[133][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11895_ (.D(_00591_),
    .CLK(net456),
    .Q(\u_cpu.rf_ram.memory[132][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11896_ (.D(_00592_),
    .CLK(net459),
    .Q(\u_cpu.rf_ram.memory[132][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11897_ (.D(_00593_),
    .CLK(net470),
    .Q(\u_cpu.rf_ram.memory[132][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11898_ (.D(_00594_),
    .CLK(net471),
    .Q(\u_cpu.rf_ram.memory[132][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11899_ (.D(_00595_),
    .CLK(net471),
    .Q(\u_cpu.rf_ram.memory[132][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11900_ (.D(_00596_),
    .CLK(net468),
    .Q(\u_cpu.rf_ram.memory[132][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11901_ (.D(_00597_),
    .CLK(net469),
    .Q(\u_cpu.rf_ram.memory[132][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11902_ (.D(_00598_),
    .CLK(net459),
    .Q(\u_cpu.rf_ram.memory[132][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11903_ (.D(_00599_),
    .CLK(net457),
    .Q(\u_cpu.rf_ram.memory[131][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11904_ (.D(_00600_),
    .CLK(net458),
    .Q(\u_cpu.rf_ram.memory[131][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11905_ (.D(_00601_),
    .CLK(net471),
    .Q(\u_cpu.rf_ram.memory[131][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11906_ (.D(_00602_),
    .CLK(net471),
    .Q(\u_cpu.rf_ram.memory[131][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11907_ (.D(_00603_),
    .CLK(net463),
    .Q(\u_cpu.rf_ram.memory[131][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11908_ (.D(_00604_),
    .CLK(net461),
    .Q(\u_cpu.rf_ram.memory[131][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11909_ (.D(_00605_),
    .CLK(net462),
    .Q(\u_cpu.rf_ram.memory[131][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11910_ (.D(_00606_),
    .CLK(net457),
    .Q(\u_cpu.rf_ram.memory[131][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11911_ (.D(_00607_),
    .CLK(net457),
    .Q(\u_cpu.rf_ram.memory[130][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11912_ (.D(_00608_),
    .CLK(net458),
    .Q(\u_cpu.rf_ram.memory[130][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11913_ (.D(_00609_),
    .CLK(net469),
    .Q(\u_cpu.rf_ram.memory[130][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11914_ (.D(_00610_),
    .CLK(net469),
    .Q(\u_cpu.rf_ram.memory[130][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11915_ (.D(_00611_),
    .CLK(net463),
    .Q(\u_cpu.rf_ram.memory[130][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11916_ (.D(_00612_),
    .CLK(net454),
    .Q(\u_cpu.rf_ram.memory[130][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11917_ (.D(_00613_),
    .CLK(net458),
    .Q(\u_cpu.rf_ram.memory[130][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11918_ (.D(_00614_),
    .CLK(net457),
    .Q(\u_cpu.rf_ram.memory[130][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11919_ (.D(_00615_),
    .CLK(net144),
    .Q(\u_cpu.rf_ram.memory[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11920_ (.D(_00616_),
    .CLK(net150),
    .Q(\u_cpu.rf_ram.memory[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11921_ (.D(_00617_),
    .CLK(net150),
    .Q(\u_cpu.rf_ram.memory[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11922_ (.D(_00618_),
    .CLK(net153),
    .Q(\u_cpu.rf_ram.memory[12][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11923_ (.D(_00619_),
    .CLK(net153),
    .Q(\u_cpu.rf_ram.memory[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11924_ (.D(_00620_),
    .CLK(net146),
    .Q(\u_cpu.rf_ram.memory[12][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11925_ (.D(_00621_),
    .CLK(net236),
    .Q(\u_cpu.rf_ram.memory[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11926_ (.D(_00622_),
    .CLK(net237),
    .Q(\u_cpu.rf_ram.memory[12][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11927_ (.D(_00623_),
    .CLK(net419),
    .Q(\u_cpu.rf_ram.memory[22][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11928_ (.D(_00624_),
    .CLK(net333),
    .Q(\u_cpu.rf_ram.memory[22][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11929_ (.D(_00625_),
    .CLK(net419),
    .Q(\u_cpu.rf_ram.memory[22][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11930_ (.D(_00626_),
    .CLK(net419),
    .Q(\u_cpu.rf_ram.memory[22][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11931_ (.D(_00627_),
    .CLK(net419),
    .Q(\u_cpu.rf_ram.memory[22][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11932_ (.D(_00628_),
    .CLK(net333),
    .Q(\u_cpu.rf_ram.memory[22][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11933_ (.D(_00629_),
    .CLK(net419),
    .Q(\u_cpu.rf_ram.memory[22][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11934_ (.D(_00630_),
    .CLK(net333),
    .Q(\u_cpu.rf_ram.memory[22][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11935_ (.D(_00631_),
    .CLK(net454),
    .Q(\u_cpu.rf_ram.memory[128][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11936_ (.D(_00632_),
    .CLK(net462),
    .Q(\u_cpu.rf_ram.memory[128][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11937_ (.D(_00633_),
    .CLK(net463),
    .Q(\u_cpu.rf_ram.memory[128][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11938_ (.D(_00634_),
    .CLK(net463),
    .Q(\u_cpu.rf_ram.memory[128][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11939_ (.D(_00635_),
    .CLK(net464),
    .Q(\u_cpu.rf_ram.memory[128][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11940_ (.D(_00636_),
    .CLK(net462),
    .Q(\u_cpu.rf_ram.memory[128][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11941_ (.D(_00637_),
    .CLK(net462),
    .Q(\u_cpu.rf_ram.memory[128][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11942_ (.D(_00638_),
    .CLK(net454),
    .Q(\u_cpu.rf_ram.memory[128][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11943_ (.D(_00639_),
    .CLK(net461),
    .Q(\u_cpu.rf_ram.memory[127][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11944_ (.D(_00640_),
    .CLK(net461),
    .Q(\u_cpu.rf_ram.memory[127][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11945_ (.D(_00641_),
    .CLK(net444),
    .Q(\u_cpu.rf_ram.memory[127][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11946_ (.D(_00642_),
    .CLK(net444),
    .Q(\u_cpu.rf_ram.memory[127][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11947_ (.D(_00643_),
    .CLK(net444),
    .Q(\u_cpu.rf_ram.memory[127][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11948_ (.D(_00644_),
    .CLK(net461),
    .Q(\u_cpu.rf_ram.memory[127][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11949_ (.D(_00645_),
    .CLK(net461),
    .Q(\u_cpu.rf_ram.memory[127][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11950_ (.D(_00646_),
    .CLK(net451),
    .Q(\u_cpu.rf_ram.memory[127][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11951_ (.D(_00647_),
    .CLK(net453),
    .Q(\u_cpu.rf_ram.memory[126][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11952_ (.D(_00648_),
    .CLK(net453),
    .Q(\u_cpu.rf_ram.memory[126][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11953_ (.D(_00649_),
    .CLK(net440),
    .Q(\u_cpu.rf_ram.memory[126][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11954_ (.D(_00650_),
    .CLK(net440),
    .Q(\u_cpu.rf_ram.memory[126][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11955_ (.D(_00651_),
    .CLK(net440),
    .Q(\u_cpu.rf_ram.memory[126][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11956_ (.D(_00652_),
    .CLK(net453),
    .Q(\u_cpu.rf_ram.memory[126][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11957_ (.D(_00653_),
    .CLK(net441),
    .Q(\u_cpu.rf_ram.memory[126][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11958_ (.D(_00654_),
    .CLK(net451),
    .Q(\u_cpu.rf_ram.memory[126][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11959_ (.D(_00655_),
    .CLK(net465),
    .Q(\u_cpu.rf_ram.memory[125][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11960_ (.D(_00656_),
    .CLK(net465),
    .Q(\u_cpu.rf_ram.memory[125][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11961_ (.D(_00657_),
    .CLK(net445),
    .Q(\u_cpu.rf_ram.memory[125][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11962_ (.D(_00658_),
    .CLK(net445),
    .Q(\u_cpu.rf_ram.memory[125][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11963_ (.D(_00659_),
    .CLK(net445),
    .Q(\u_cpu.rf_ram.memory[125][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11964_ (.D(_00660_),
    .CLK(net465),
    .Q(\u_cpu.rf_ram.memory[125][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11965_ (.D(_00661_),
    .CLK(net465),
    .Q(\u_cpu.rf_ram.memory[125][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11966_ (.D(_00662_),
    .CLK(net453),
    .Q(\u_cpu.rf_ram.memory[125][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11967_ (.D(_00663_),
    .CLK(net464),
    .Q(\u_cpu.rf_ram.memory[124][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11968_ (.D(_00664_),
    .CLK(net463),
    .Q(\u_cpu.rf_ram.memory[124][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11969_ (.D(_00665_),
    .CLK(net446),
    .Q(\u_cpu.rf_ram.memory[124][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11970_ (.D(_00666_),
    .CLK(net445),
    .Q(\u_cpu.rf_ram.memory[124][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11971_ (.D(_00667_),
    .CLK(net445),
    .Q(\u_cpu.rf_ram.memory[124][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11972_ (.D(_00668_),
    .CLK(net465),
    .Q(\u_cpu.rf_ram.memory[124][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11973_ (.D(_00669_),
    .CLK(net446),
    .Q(\u_cpu.rf_ram.memory[124][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11974_ (.D(_00670_),
    .CLK(net453),
    .Q(\u_cpu.rf_ram.memory[124][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11975_ (.D(_00015_),
    .CLK(net263),
    .Q(\u_cpu.rf_ram_if.rdata1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11976_ (.D(_00016_),
    .CLK(net265),
    .Q(\u_cpu.rf_ram_if.rdata1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11977_ (.D(_00017_),
    .CLK(net265),
    .Q(\u_cpu.rf_ram_if.rdata1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11978_ (.D(_00018_),
    .CLK(net265),
    .Q(\u_cpu.rf_ram_if.rdata1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11979_ (.D(_00019_),
    .CLK(net265),
    .Q(\u_cpu.rf_ram_if.rdata1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11980_ (.D(_00020_),
    .CLK(net254),
    .Q(\u_cpu.rf_ram_if.rdata1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11981_ (.D(_00671_),
    .CLK(net410),
    .Q(\u_cpu.rf_ram.memory[123][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11982_ (.D(_00672_),
    .CLK(net411),
    .Q(\u_cpu.rf_ram.memory[123][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11983_ (.D(_00673_),
    .CLK(net410),
    .Q(\u_cpu.rf_ram.memory[123][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11984_ (.D(_00674_),
    .CLK(net438),
    .Q(\u_cpu.rf_ram.memory[123][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11985_ (.D(_00675_),
    .CLK(net438),
    .Q(\u_cpu.rf_ram.memory[123][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11986_ (.D(_00676_),
    .CLK(net439),
    .Q(\u_cpu.rf_ram.memory[123][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11987_ (.D(_00677_),
    .CLK(net439),
    .Q(\u_cpu.rf_ram.memory[123][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11988_ (.D(_00678_),
    .CLK(net439),
    .Q(\u_cpu.rf_ram.memory[123][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11989_ (.D(_00008_),
    .CLK(net263),
    .Q(\u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11990_ (.D(_00009_),
    .CLK(net263),
    .Q(\u_cpu.rf_ram_if.rdata0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11991_ (.D(_00010_),
    .CLK(net257),
    .Q(\u_cpu.rf_ram_if.rdata0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11992_ (.D(_00011_),
    .CLK(net259),
    .Q(\u_cpu.rf_ram_if.rdata0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11993_ (.D(_00012_),
    .CLK(net259),
    .Q(\u_cpu.rf_ram_if.rdata0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11994_ (.D(_00013_),
    .CLK(net259),
    .Q(\u_cpu.rf_ram_if.rdata0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11995_ (.D(_00014_),
    .CLK(net257),
    .Q(\u_cpu.rf_ram_if.rdata0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11996_ (.D(_00679_),
    .CLK(net400),
    .Q(\u_cpu.rf_ram.memory[38][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11997_ (.D(_00680_),
    .CLK(net400),
    .Q(\u_cpu.rf_ram.memory[38][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11998_ (.D(_00681_),
    .CLK(net400),
    .Q(\u_cpu.rf_ram.memory[38][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11999_ (.D(_00682_),
    .CLK(net401),
    .Q(\u_cpu.rf_ram.memory[38][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12000_ (.D(_00683_),
    .CLK(net401),
    .Q(\u_cpu.rf_ram.memory[38][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12001_ (.D(_00684_),
    .CLK(net415),
    .Q(\u_cpu.rf_ram.memory[38][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12002_ (.D(_00685_),
    .CLK(net415),
    .Q(\u_cpu.rf_ram.memory[38][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12003_ (.D(_00686_),
    .CLK(net415),
    .Q(\u_cpu.rf_ram.memory[38][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12004_ (.D(_00687_),
    .CLK(net408),
    .Q(\u_cpu.rf_ram.memory[37][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12005_ (.D(_00688_),
    .CLK(net408),
    .Q(\u_cpu.rf_ram.memory[37][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12006_ (.D(_00689_),
    .CLK(net409),
    .Q(\u_cpu.rf_ram.memory[37][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12007_ (.D(_00690_),
    .CLK(net409),
    .Q(\u_cpu.rf_ram.memory[37][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12008_ (.D(_00691_),
    .CLK(net409),
    .Q(\u_cpu.rf_ram.memory[37][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12009_ (.D(_00692_),
    .CLK(net425),
    .Q(\u_cpu.rf_ram.memory[37][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12010_ (.D(_00693_),
    .CLK(net425),
    .Q(\u_cpu.rf_ram.memory[37][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12011_ (.D(_00694_),
    .CLK(net425),
    .Q(\u_cpu.rf_ram.memory[37][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12012_ (.D(_00695_),
    .CLK(net411),
    .Q(\u_cpu.rf_ram.memory[36][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12013_ (.D(_00696_),
    .CLK(net411),
    .Q(\u_cpu.rf_ram.memory[36][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12014_ (.D(_00697_),
    .CLK(net411),
    .Q(\u_cpu.rf_ram.memory[36][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12015_ (.D(_00698_),
    .CLK(net439),
    .Q(\u_cpu.rf_ram.memory[36][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12016_ (.D(_00699_),
    .CLK(net439),
    .Q(\u_cpu.rf_ram.memory[36][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12017_ (.D(_00700_),
    .CLK(net450),
    .Q(\u_cpu.rf_ram.memory[36][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12018_ (.D(_00701_),
    .CLK(net450),
    .Q(\u_cpu.rf_ram.memory[36][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12019_ (.D(_00702_),
    .CLK(net428),
    .Q(\u_cpu.rf_ram.memory[36][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12020_ (.D(_00703_),
    .CLK(net379),
    .Q(\u_cpu.cpu.state.stage_two_req ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12021_ (.D(_00704_),
    .CLK(net481),
    .Q(\u_cpu.cpu.state.o_cnt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12022_ (.D(_00705_),
    .CLK(net482),
    .Q(\u_cpu.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12023_ (.D(_00706_),
    .CLK(net495),
    .Q(\u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12024_ (.D(_00707_),
    .CLK(net482),
    .Q(\u_cpu.cpu.state.o_cnt_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12025_ (.D(_00708_),
    .CLK(net490),
    .Q(\u_cpu.cpu.state.o_cnt_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12026_ (.D(_00709_),
    .CLK(net490),
    .Q(\u_cpu.cpu.state.o_cnt_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12027_ (.D(_00710_),
    .CLK(net492),
    .Q(\u_cpu.cpu.state.o_cnt_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12028_ (.D(_00711_),
    .CLK(net320),
    .Q(\u_cpu.rf_ram.memory[91][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12029_ (.D(_00712_),
    .CLK(net313),
    .Q(\u_cpu.rf_ram.memory[91][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12030_ (.D(_00713_),
    .CLK(net312),
    .Q(\u_cpu.rf_ram.memory[91][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12031_ (.D(_00714_),
    .CLK(net312),
    .Q(\u_cpu.rf_ram.memory[91][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12032_ (.D(_00715_),
    .CLK(net312),
    .Q(\u_cpu.rf_ram.memory[91][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12033_ (.D(_00716_),
    .CLK(net319),
    .Q(\u_cpu.rf_ram.memory[91][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12034_ (.D(_00717_),
    .CLK(net319),
    .Q(\u_cpu.rf_ram.memory[91][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12035_ (.D(_00718_),
    .CLK(net313),
    .Q(\u_cpu.rf_ram.memory[91][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12036_ (.D(_00719_),
    .CLK(net284),
    .Q(\u_cpu.rf_ram.memory[90][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12037_ (.D(_00720_),
    .CLK(net284),
    .Q(\u_cpu.rf_ram.memory[90][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12038_ (.D(_00721_),
    .CLK(net285),
    .Q(\u_cpu.rf_ram.memory[90][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12039_ (.D(_00722_),
    .CLK(net285),
    .Q(\u_cpu.rf_ram.memory[90][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12040_ (.D(_00723_),
    .CLK(net285),
    .Q(\u_cpu.rf_ram.memory[90][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12041_ (.D(_00724_),
    .CLK(net308),
    .Q(\u_cpu.rf_ram.memory[90][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12042_ (.D(_00725_),
    .CLK(net308),
    .Q(\u_cpu.rf_ram.memory[90][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12043_ (.D(_00726_),
    .CLK(net308),
    .Q(\u_cpu.rf_ram.memory[90][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12044_ (.D(_00727_),
    .CLK(net480),
    .Q(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12045_ (.D(_00728_),
    .CLK(net495),
    .Q(\u_cpu.cpu.mem_if.signbit ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12046_ (.D(_00729_),
    .CLK(net495),
    .Q(\u_cpu.cpu.ctrl.i_jump ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12047_ (.D(_00730_),
    .CLK(net500),
    .Q(\u_cpu.cpu.bufreg2.i_cnt_done ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12048_ (.D(_00731_),
    .CLK(net379),
    .Q(\u_cpu.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12049_ (.D(_00732_),
    .CLK(net271),
    .Q(\u_cpu.rf_ram.memory[92][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12050_ (.D(_00733_),
    .CLK(net270),
    .Q(\u_cpu.rf_ram.memory[92][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12051_ (.D(_00734_),
    .CLK(net270),
    .Q(\u_cpu.rf_ram.memory[92][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12052_ (.D(_00735_),
    .CLK(net270),
    .Q(\u_cpu.rf_ram.memory[92][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12053_ (.D(_00736_),
    .CLK(net270),
    .Q(\u_cpu.rf_ram.memory[92][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12054_ (.D(_00737_),
    .CLK(net270),
    .Q(\u_cpu.rf_ram.memory[92][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12055_ (.D(_00738_),
    .CLK(net271),
    .Q(\u_cpu.rf_ram.memory[92][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12056_ (.D(_00739_),
    .CLK(net271),
    .Q(\u_cpu.rf_ram.memory[92][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12057_ (.D(_00740_),
    .CLK(net308),
    .Q(\u_cpu.rf_ram.memory[35][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12058_ (.D(_00741_),
    .CLK(net307),
    .Q(\u_cpu.rf_ram.memory[35][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12059_ (.D(_00742_),
    .CLK(net307),
    .Q(\u_cpu.rf_ram.memory[35][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12060_ (.D(_00743_),
    .CLK(net307),
    .Q(\u_cpu.rf_ram.memory[35][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12061_ (.D(_00744_),
    .CLK(net307),
    .Q(\u_cpu.rf_ram.memory[35][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12062_ (.D(_00745_),
    .CLK(net285),
    .Q(\u_cpu.rf_ram.memory[35][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12063_ (.D(_00746_),
    .CLK(net307),
    .Q(\u_cpu.rf_ram.memory[35][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12064_ (.D(_00747_),
    .CLK(net289),
    .Q(\u_cpu.rf_ram.memory[35][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12065_ (.D(_00748_),
    .CLK(net284),
    .Q(\u_cpu.rf_ram.memory[34][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12066_ (.D(_00749_),
    .CLK(net282),
    .Q(\u_cpu.rf_ram.memory[34][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12067_ (.D(_00750_),
    .CLK(net282),
    .Q(\u_cpu.rf_ram.memory[34][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12068_ (.D(_00751_),
    .CLK(net282),
    .Q(\u_cpu.rf_ram.memory[34][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12069_ (.D(_00752_),
    .CLK(net282),
    .Q(\u_cpu.rf_ram.memory[34][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12070_ (.D(_00753_),
    .CLK(net282),
    .Q(\u_cpu.rf_ram.memory[34][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12071_ (.D(_00754_),
    .CLK(net283),
    .Q(\u_cpu.rf_ram.memory[34][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12072_ (.D(_00755_),
    .CLK(net284),
    .Q(\u_cpu.rf_ram.memory[34][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12073_ (.D(_00756_),
    .CLK(net310),
    .Q(\u_cpu.rf_ram.memory[117][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12074_ (.D(_00757_),
    .CLK(net312),
    .Q(\u_cpu.rf_ram.memory[117][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12075_ (.D(_00758_),
    .CLK(net318),
    .Q(\u_cpu.rf_ram.memory[117][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12076_ (.D(_00759_),
    .CLK(net318),
    .Q(\u_cpu.rf_ram.memory[117][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12077_ (.D(_00760_),
    .CLK(net310),
    .Q(\u_cpu.rf_ram.memory[117][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12078_ (.D(_00761_),
    .CLK(net319),
    .Q(\u_cpu.rf_ram.memory[117][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12079_ (.D(_00762_),
    .CLK(net319),
    .Q(\u_cpu.rf_ram.memory[117][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12080_ (.D(_00763_),
    .CLK(net312),
    .Q(\u_cpu.rf_ram.memory[117][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12081_ (.D(_00764_),
    .CLK(net410),
    .Q(\u_cpu.rf_ram.memory[120][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12082_ (.D(_00765_),
    .CLK(net436),
    .Q(\u_cpu.rf_ram.memory[120][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12083_ (.D(_00766_),
    .CLK(net448),
    .Q(\u_cpu.rf_ram.memory[120][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12084_ (.D(_00767_),
    .CLK(net437),
    .Q(\u_cpu.rf_ram.memory[120][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12085_ (.D(_00768_),
    .CLK(net443),
    .Q(\u_cpu.rf_ram.memory[120][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12086_ (.D(_00769_),
    .CLK(net443),
    .Q(\u_cpu.rf_ram.memory[120][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12087_ (.D(_00770_),
    .CLK(net443),
    .Q(\u_cpu.rf_ram.memory[120][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12088_ (.D(_00771_),
    .CLK(net438),
    .Q(\u_cpu.rf_ram.memory[120][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12089_ (.D(_00772_),
    .CLK(net401),
    .Q(\u_cpu.rf_ram.memory[118][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12090_ (.D(_00773_),
    .CLK(net401),
    .Q(\u_cpu.rf_ram.memory[118][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12091_ (.D(_00774_),
    .CLK(net403),
    .Q(\u_cpu.rf_ram.memory[118][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12092_ (.D(_00775_),
    .CLK(net404),
    .Q(\u_cpu.rf_ram.memory[118][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12093_ (.D(_00776_),
    .CLK(net404),
    .Q(\u_cpu.rf_ram.memory[118][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12094_ (.D(_00777_),
    .CLK(net408),
    .Q(\u_cpu.rf_ram.memory[118][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12095_ (.D(_00778_),
    .CLK(net408),
    .Q(\u_cpu.rf_ram.memory[118][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12096_ (.D(_00779_),
    .CLK(net408),
    .Q(\u_cpu.rf_ram.memory[118][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12097_ (.D(_00780_),
    .CLK(net410),
    .Q(\u_cpu.rf_ram.memory[121][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12098_ (.D(_00781_),
    .CLK(net405),
    .Q(\u_cpu.rf_ram.memory[121][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12099_ (.D(_00782_),
    .CLK(net448),
    .Q(\u_cpu.rf_ram.memory[121][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12100_ (.D(_00783_),
    .CLK(net437),
    .Q(\u_cpu.rf_ram.memory[121][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12101_ (.D(_00784_),
    .CLK(net443),
    .Q(\u_cpu.rf_ram.memory[121][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12102_ (.D(_00785_),
    .CLK(net444),
    .Q(\u_cpu.rf_ram.memory[121][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12103_ (.D(_00786_),
    .CLK(net443),
    .Q(\u_cpu.rf_ram.memory[121][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12104_ (.D(_00787_),
    .CLK(net441),
    .Q(\u_cpu.rf_ram.memory[121][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12105_ (.D(_00788_),
    .CLK(net125),
    .Q(\u_cpu.rf_ram.memory[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12106_ (.D(_00789_),
    .CLK(net125),
    .Q(\u_cpu.rf_ram.memory[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12107_ (.D(_00790_),
    .CLK(net118),
    .Q(\u_cpu.rf_ram.memory[8][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12108_ (.D(_00791_),
    .CLK(net117),
    .Q(\u_cpu.rf_ram.memory[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12109_ (.D(_00792_),
    .CLK(net128),
    .Q(\u_cpu.rf_ram.memory[8][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12110_ (.D(_00793_),
    .CLK(net127),
    .Q(\u_cpu.rf_ram.memory[8][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12111_ (.D(_00794_),
    .CLK(net143),
    .Q(\u_cpu.rf_ram.memory[8][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12112_ (.D(_00795_),
    .CLK(net137),
    .Q(\u_cpu.rf_ram.memory[8][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12113_ (.D(_00796_),
    .CLK(net125),
    .Q(\u_cpu.rf_ram.memory[11][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12114_ (.D(_00797_),
    .CLK(net118),
    .Q(\u_cpu.rf_ram.memory[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12115_ (.D(_00798_),
    .CLK(net116),
    .Q(\u_cpu.rf_ram.memory[11][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12116_ (.D(_00799_),
    .CLK(net116),
    .Q(\u_cpu.rf_ram.memory[11][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12117_ (.D(_00800_),
    .CLK(net128),
    .Q(\u_cpu.rf_ram.memory[11][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12118_ (.D(_00801_),
    .CLK(net127),
    .Q(\u_cpu.rf_ram.memory[11][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12119_ (.D(_00802_),
    .CLK(net143),
    .Q(\u_cpu.rf_ram.memory[11][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12120_ (.D(_00803_),
    .CLK(net137),
    .Q(\u_cpu.rf_ram.memory[11][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12121_ (.D(_00804_),
    .CLK(net405),
    .Q(\u_cpu.rf_ram.memory[112][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12122_ (.D(_00805_),
    .CLK(net406),
    .Q(\u_cpu.rf_ram.memory[112][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12123_ (.D(_00806_),
    .CLK(net406),
    .Q(\u_cpu.rf_ram.memory[112][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12124_ (.D(_00807_),
    .CLK(net406),
    .Q(\u_cpu.rf_ram.memory[112][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12125_ (.D(_00808_),
    .CLK(net406),
    .Q(\u_cpu.rf_ram.memory[112][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12126_ (.D(_00809_),
    .CLK(net405),
    .Q(\u_cpu.rf_ram.memory[112][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12127_ (.D(_00810_),
    .CLK(net407),
    .Q(\u_cpu.rf_ram.memory[112][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12128_ (.D(_00811_),
    .CLK(net405),
    .Q(\u_cpu.rf_ram.memory[112][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12129_ (.D(_00812_),
    .CLK(net410),
    .Q(\u_cpu.rf_ram.memory[122][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12130_ (.D(_00813_),
    .CLK(net405),
    .Q(\u_cpu.rf_ram.memory[122][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12131_ (.D(_00814_),
    .CLK(net436),
    .Q(\u_cpu.rf_ram.memory[122][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12132_ (.D(_00815_),
    .CLK(net436),
    .Q(\u_cpu.rf_ram.memory[122][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12133_ (.D(_00816_),
    .CLK(net436),
    .Q(\u_cpu.rf_ram.memory[122][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12134_ (.D(_00817_),
    .CLK(net438),
    .Q(\u_cpu.rf_ram.memory[122][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12135_ (.D(_00818_),
    .CLK(net436),
    .Q(\u_cpu.rf_ram.memory[122][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12136_ (.D(_00819_),
    .CLK(net438),
    .Q(\u_cpu.rf_ram.memory[122][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12137_ (.D(_00820_),
    .CLK(net403),
    .Q(\u_cpu.rf_ram.memory[115][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12138_ (.D(_00821_),
    .CLK(net403),
    .Q(\u_cpu.rf_ram.memory[115][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12139_ (.D(_00822_),
    .CLK(net398),
    .Q(\u_cpu.rf_ram.memory[115][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12140_ (.D(_00823_),
    .CLK(net396),
    .Q(\u_cpu.rf_ram.memory[115][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12141_ (.D(_00824_),
    .CLK(net396),
    .Q(\u_cpu.rf_ram.memory[115][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12142_ (.D(_00825_),
    .CLK(net317),
    .Q(\u_cpu.rf_ram.memory[115][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12143_ (.D(_00826_),
    .CLK(net396),
    .Q(\u_cpu.rf_ram.memory[115][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12144_ (.D(_00827_),
    .CLK(net398),
    .Q(\u_cpu.rf_ram.memory[115][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12145_ (.D(_00828_),
    .CLK(net397),
    .Q(\u_cpu.rf_ram.memory[116][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12146_ (.D(_00829_),
    .CLK(net397),
    .Q(\u_cpu.rf_ram.memory[116][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12147_ (.D(_00830_),
    .CLK(net317),
    .Q(\u_cpu.rf_ram.memory[116][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12148_ (.D(_00831_),
    .CLK(net317),
    .Q(\u_cpu.rf_ram.memory[116][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12149_ (.D(_00832_),
    .CLK(net317),
    .Q(\u_cpu.rf_ram.memory[116][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12150_ (.D(_00833_),
    .CLK(net397),
    .Q(\u_cpu.rf_ram.memory[116][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12151_ (.D(_00834_),
    .CLK(net401),
    .Q(\u_cpu.rf_ram.memory[116][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12152_ (.D(_00835_),
    .CLK(net398),
    .Q(\u_cpu.rf_ram.memory[116][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12153_ (.D(_00836_),
    .CLK(net310),
    .Q(\u_cpu.rf_ram.memory[33][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12154_ (.D(_00837_),
    .CLK(net309),
    .Q(\u_cpu.rf_ram.memory[33][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12155_ (.D(_00838_),
    .CLK(net309),
    .Q(\u_cpu.rf_ram.memory[33][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12156_ (.D(_00839_),
    .CLK(net309),
    .Q(\u_cpu.rf_ram.memory[33][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12157_ (.D(_00840_),
    .CLK(net309),
    .Q(\u_cpu.rf_ram.memory[33][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12158_ (.D(_00841_),
    .CLK(net309),
    .Q(\u_cpu.rf_ram.memory[33][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12159_ (.D(_00842_),
    .CLK(net310),
    .Q(\u_cpu.rf_ram.memory[33][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12160_ (.D(_00843_),
    .CLK(net311),
    .Q(\u_cpu.rf_ram.memory[33][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12161_ (.D(_00844_),
    .CLK(net497),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12162_ (.D(_00845_),
    .CLK(net497),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12163_ (.D(_00846_),
    .CLK(net498),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12164_ (.D(_00847_),
    .CLK(net390),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12165_ (.D(_00848_),
    .CLK(net390),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12166_ (.D(_00849_),
    .CLK(net391),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12167_ (.D(_00850_),
    .CLK(net389),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12168_ (.D(_00851_),
    .CLK(net387),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12169_ (.D(_00852_),
    .CLK(net385),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12170_ (.D(_00853_),
    .CLK(net383),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12171_ (.D(_00854_),
    .CLK(net386),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12172_ (.D(_00855_),
    .CLK(net386),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12173_ (.D(_00856_),
    .CLK(net386),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12174_ (.D(_00857_),
    .CLK(net363),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12175_ (.D(_00858_),
    .CLK(net386),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12176_ (.D(_00859_),
    .CLK(net387),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12177_ (.D(_00860_),
    .CLK(net387),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12178_ (.D(_00861_),
    .CLK(net386),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12179_ (.D(_00862_),
    .CLK(net387),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12180_ (.D(_00863_),
    .CLK(net388),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12181_ (.D(_00864_),
    .CLK(net389),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12182_ (.D(_00865_),
    .CLK(net389),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12183_ (.D(_00866_),
    .CLK(net389),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12184_ (.D(_00867_),
    .CLK(net389),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12185_ (.D(_00868_),
    .CLK(net390),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12186_ (.D(_00869_),
    .CLK(net497),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12187_ (.D(_00870_),
    .CLK(net497),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12188_ (.D(_00871_),
    .CLK(net390),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12189_ (.D(_00872_),
    .CLK(net497),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12190_ (.D(_00873_),
    .CLK(net498),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12191_ (.D(_00874_),
    .CLK(net498),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12192_ (.D(_00875_),
    .CLK(net498),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12193_ (.D(_00876_),
    .CLK(net403),
    .Q(\u_cpu.rf_ram.memory[113][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12194_ (.D(_00877_),
    .CLK(net403),
    .Q(\u_cpu.rf_ram.memory[113][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12195_ (.D(_00878_),
    .CLK(net398),
    .Q(\u_cpu.rf_ram.memory[113][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12196_ (.D(_00879_),
    .CLK(net396),
    .Q(\u_cpu.rf_ram.memory[113][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12197_ (.D(_00880_),
    .CLK(net396),
    .Q(\u_cpu.rf_ram.memory[113][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12198_ (.D(_00881_),
    .CLK(net397),
    .Q(\u_cpu.rf_ram.memory[113][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12199_ (.D(_00882_),
    .CLK(net398),
    .Q(\u_cpu.rf_ram.memory[113][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12200_ (.D(_00883_),
    .CLK(net399),
    .Q(\u_cpu.rf_ram.memory[113][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12201_ (.D(_00884_),
    .CLK(net384),
    .Q(\u_cpu.cpu.decode.opcode[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12202_ (.D(_00885_),
    .CLK(net360),
    .Q(\u_cpu.cpu.decode.opcode[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12203_ (.D(_00886_),
    .CLK(net384),
    .Q(\u_cpu.cpu.decode.opcode[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12204_ (.D(_00887_),
    .CLK(net362),
    .Q(\u_arbiter.i_wb_cpu_dbus_we ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12205_ (.D(_00888_),
    .CLK(net384),
    .Q(\u_cpu.cpu.branch_op ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12206_ (.D(_00889_),
    .CLK(net383),
    .Q(\u_cpu.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12207_ (.D(_00890_),
    .CLK(net385),
    .Q(\u_cpu.cpu.decode.co_mem_word ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12208_ (.D(_00891_),
    .CLK(net384),
    .Q(\u_cpu.cpu.csr_d_sel ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12209_ (.D(_00892_),
    .CLK(net373),
    .Q(\u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12210_ (.D(_00893_),
    .CLK(net352),
    .Q(\u_cpu.cpu.decode.op21 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12211_ (.D(_00894_),
    .CLK(net353),
    .Q(\u_cpu.cpu.decode.op22 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12212_ (.D(_00895_),
    .CLK(net318),
    .Q(\u_cpu.rf_ram.memory[114][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12213_ (.D(_00896_),
    .CLK(net318),
    .Q(\u_cpu.rf_ram.memory[114][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12214_ (.D(_00897_),
    .CLK(net316),
    .Q(\u_cpu.rf_ram.memory[114][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12215_ (.D(_00898_),
    .CLK(net316),
    .Q(\u_cpu.rf_ram.memory[114][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12216_ (.D(_00899_),
    .CLK(net316),
    .Q(\u_cpu.rf_ram.memory[114][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12217_ (.D(_00900_),
    .CLK(net316),
    .Q(\u_cpu.rf_ram.memory[114][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12218_ (.D(_00901_),
    .CLK(net316),
    .Q(\u_cpu.rf_ram.memory[114][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12219_ (.D(_00902_),
    .CLK(net318),
    .Q(\u_cpu.rf_ram.memory[114][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12220_ (.D(_00903_),
    .CLK(net353),
    .Q(\u_cpu.cpu.decode.op26 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12221_ (.D(_00904_),
    .CLK(net350),
    .Q(\u_cpu.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12222_ (.D(_00905_),
    .CLK(net351),
    .Q(\u_cpu.cpu.immdec.imm24_20[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12223_ (.D(_00906_),
    .CLK(net343),
    .Q(\u_cpu.cpu.immdec.imm24_20[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12224_ (.D(_00907_),
    .CLK(net343),
    .Q(\u_cpu.cpu.immdec.imm24_20[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12225_ (.D(_00908_),
    .CLK(net359),
    .Q(\u_cpu.cpu.immdec.imm24_20[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12226_ (.D(_00909_),
    .CLK(net362),
    .Q(\u_cpu.cpu.immdec.imm30_25[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12227_ (.D(_00910_),
    .CLK(net360),
    .Q(\u_cpu.cpu.immdec.imm30_25[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12228_ (.D(_00911_),
    .CLK(net360),
    .Q(\u_cpu.cpu.immdec.imm30_25[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12229_ (.D(_00912_),
    .CLK(net361),
    .Q(\u_cpu.cpu.immdec.imm30_25[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12230_ (.D(_00913_),
    .CLK(net361),
    .Q(\u_cpu.cpu.immdec.imm30_25[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12231_ (.D(_00914_),
    .CLK(net383),
    .Q(\u_cpu.cpu.immdec.imm30_25[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12232_ (.D(_00915_),
    .CLK(net360),
    .Q(\u_cpu.cpu.immdec.imm7 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12233_ (.D(_00916_),
    .CLK(net359),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12234_ (.D(_00917_),
    .CLK(net263),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12235_ (.D(_00918_),
    .CLK(net263),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12236_ (.D(_00919_),
    .CLK(net264),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12237_ (.D(_00920_),
    .CLK(net359),
    .Q(\u_cpu.cpu.csr_imm ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12238_ (.D(_00921_),
    .CLK(net341),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12239_ (.D(_00922_),
    .CLK(net341),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12240_ (.D(_00923_),
    .CLK(net342),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12241_ (.D(_00924_),
    .CLK(net260),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12242_ (.D(_00925_),
    .CLK(net383),
    .Q(\u_cpu.cpu.immdec.imm31 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12243_ (.D(_00926_),
    .CLK(net480),
    .Q(\u_cpu.cpu.genblk3.csr.timer_irq_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12244_ (.D(_00927_),
    .CLK(net274),
    .Q(\u_cpu.rf_ram.memory[32][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12245_ (.D(_00928_),
    .CLK(net272),
    .Q(\u_cpu.rf_ram.memory[32][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12246_ (.D(_00929_),
    .CLK(net272),
    .Q(\u_cpu.rf_ram.memory[32][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12247_ (.D(_00930_),
    .CLK(net272),
    .Q(\u_cpu.rf_ram.memory[32][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12248_ (.D(_00931_),
    .CLK(net272),
    .Q(\u_cpu.rf_ram.memory[32][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12249_ (.D(_00932_),
    .CLK(net272),
    .Q(\u_cpu.rf_ram.memory[32][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12250_ (.D(_00933_),
    .CLK(net273),
    .Q(\u_cpu.rf_ram.memory[32][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12251_ (.D(_00934_),
    .CLK(net274),
    .Q(\u_cpu.rf_ram.memory[32][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12252_ (.D(_00935_),
    .CLK(net93),
    .Q(\u_cpu.rf_ram.memory[31][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12253_ (.D(_00936_),
    .CLK(net93),
    .Q(\u_cpu.rf_ram.memory[31][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12254_ (.D(_00937_),
    .CLK(net97),
    .Q(\u_cpu.rf_ram.memory[31][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12255_ (.D(_00938_),
    .CLK(net103),
    .Q(\u_cpu.rf_ram.memory[31][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12256_ (.D(_00939_),
    .CLK(net93),
    .Q(\u_cpu.rf_ram.memory[31][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12257_ (.D(_00940_),
    .CLK(net81),
    .Q(\u_cpu.rf_ram.memory[31][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12258_ (.D(_00941_),
    .CLK(net79),
    .Q(\u_cpu.rf_ram.memory[31][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12259_ (.D(_00942_),
    .CLK(net90),
    .Q(\u_cpu.rf_ram.memory[31][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12260_ (.D(_00943_),
    .CLK(net391),
    .Q(\u_cpu.cpu.alu.cmp_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12261_ (.D(_00944_),
    .CLK(net491),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12262_ (.D(_00945_),
    .CLK(net491),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12263_ (.D(_00946_),
    .CLK(net513),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12264_ (.D(_00947_),
    .CLK(net513),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12265_ (.D(_00948_),
    .CLK(net515),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12266_ (.D(_00949_),
    .CLK(net521),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12267_ (.D(_00950_),
    .CLK(net521),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12268_ (.D(_00951_),
    .CLK(net521),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12269_ (.D(_00952_),
    .CLK(net530),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12270_ (.D(_00953_),
    .CLK(net530),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12271_ (.D(_00954_),
    .CLK(net530),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12272_ (.D(_00955_),
    .CLK(net531),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12273_ (.D(_00956_),
    .CLK(net531),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12274_ (.D(_00957_),
    .CLK(net533),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12275_ (.D(_00958_),
    .CLK(net533),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12276_ (.D(_00959_),
    .CLK(net533),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12277_ (.D(_00960_),
    .CLK(net533),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12278_ (.D(_00961_),
    .CLK(net532),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12279_ (.D(_00962_),
    .CLK(net525),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12280_ (.D(_00963_),
    .CLK(net526),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12281_ (.D(_00964_),
    .CLK(net525),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12282_ (.D(_00965_),
    .CLK(net525),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12283_ (.D(_00966_),
    .CLK(net504),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12284_ (.D(_00967_),
    .CLK(net504),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12285_ (.D(_00968_),
    .CLK(net505),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12286_ (.D(_00969_),
    .CLK(net502),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12287_ (.D(_00970_),
    .CLK(net502),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12288_ (.D(_00971_),
    .CLK(net523),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12289_ (.D(_00972_),
    .CLK(net500),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12290_ (.D(_00973_),
    .CLK(net501),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12291_ (.D(_00022_),
    .CLK(net495),
    .Q(\u_cpu.cpu.bufreg.c_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12292_ (.D(_00974_),
    .CLK(net495),
    .Q(\u_cpu.cpu.bufreg.lsb[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12293_ (.D(_00975_),
    .CLK(net496),
    .Q(\u_cpu.cpu.bufreg.lsb[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12294_ (.D(_00976_),
    .CLK(net94),
    .Q(\u_cpu.rf_ram.memory[30][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12295_ (.D(_00977_),
    .CLK(net93),
    .Q(\u_cpu.rf_ram.memory[30][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12296_ (.D(_00978_),
    .CLK(net97),
    .Q(\u_cpu.rf_ram.memory[30][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12297_ (.D(_00979_),
    .CLK(net103),
    .Q(\u_cpu.rf_ram.memory[30][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12298_ (.D(_00980_),
    .CLK(net94),
    .Q(\u_cpu.rf_ram.memory[30][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12299_ (.D(_00981_),
    .CLK(net81),
    .Q(\u_cpu.rf_ram.memory[30][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12300_ (.D(_00982_),
    .CLK(net79),
    .Q(\u_cpu.rf_ram.memory[30][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12301_ (.D(_00983_),
    .CLK(net90),
    .Q(\u_cpu.rf_ram.memory[30][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12302_ (.D(_00024_),
    .CLK(net496),
    .Q(\u_cpu.cpu.ctrl.pc_plus_offset_cy_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12303_ (.D(_00023_),
    .CLK(net500),
    .Q(\u_cpu.cpu.ctrl.pc_plus_4_cy_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12304_ (.D(_00984_),
    .CLK(net500),
    .Q(\u_arbiter.i_wb_cpu_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12305_ (.D(_00985_),
    .CLK(net502),
    .Q(\u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12306_ (.D(_00986_),
    .CLK(net503),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12307_ (.D(_00987_),
    .CLK(net492),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12308_ (.D(_00988_),
    .CLK(net523),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12309_ (.D(_00989_),
    .CLK(net523),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12310_ (.D(_00990_),
    .CLK(net524),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12311_ (.D(_00991_),
    .CLK(net528),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12312_ (.D(_00992_),
    .CLK(net528),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12313_ (.D(_00993_),
    .CLK(net528),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12314_ (.D(_00994_),
    .CLK(net528),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12315_ (.D(_00995_),
    .CLK(net528),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12316_ (.D(_00996_),
    .CLK(net529),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12317_ (.D(_00997_),
    .CLK(net524),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12318_ (.D(_00998_),
    .CLK(net529),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12319_ (.D(_00999_),
    .CLK(net532),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12320_ (.D(_01000_),
    .CLK(net532),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12321_ (.D(_01001_),
    .CLK(net532),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12322_ (.D(_01002_),
    .CLK(net532),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12323_ (.D(_01003_),
    .CLK(net526),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12324_ (.D(_01004_),
    .CLK(net526),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12325_ (.D(_01005_),
    .CLK(net526),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12326_ (.D(_01006_),
    .CLK(net525),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12327_ (.D(_01007_),
    .CLK(net525),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12328_ (.D(_01008_),
    .CLK(net504),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12329_ (.D(_01009_),
    .CLK(net504),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12330_ (.D(_01010_),
    .CLK(net504),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12331_ (.D(_01011_),
    .CLK(net501),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12332_ (.D(_01012_),
    .CLK(net501),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12333_ (.D(_01013_),
    .CLK(net503),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12334_ (.D(_01014_),
    .CLK(net523),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12335_ (.D(_01015_),
    .CLK(net523),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12336_ (.D(_01016_),
    .CLK(net167),
    .Q(\u_cpu.rf_ram.memory[109][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12337_ (.D(_01017_),
    .CLK(net167),
    .Q(\u_cpu.rf_ram.memory[109][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12338_ (.D(_01018_),
    .CLK(net167),
    .Q(\u_cpu.rf_ram.memory[109][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12339_ (.D(_01019_),
    .CLK(net165),
    .Q(\u_cpu.rf_ram.memory[109][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12340_ (.D(_01020_),
    .CLK(net165),
    .Q(\u_cpu.rf_ram.memory[109][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12341_ (.D(_01021_),
    .CLK(net165),
    .Q(\u_cpu.rf_ram.memory[109][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12342_ (.D(_01022_),
    .CLK(net165),
    .Q(\u_cpu.rf_ram.memory[109][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12343_ (.D(_01023_),
    .CLK(net165),
    .Q(\u_cpu.rf_ram.memory[109][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12344_ (.D(_00021_),
    .CLK(net385),
    .Q(\u_cpu.cpu.alu.add_cy_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12345_ (.D(_01024_),
    .CLK(net112),
    .Q(\u_cpu.rf_ram.memory[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12346_ (.D(_01025_),
    .CLK(net117),
    .Q(\u_cpu.rf_ram.memory[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12347_ (.D(_01026_),
    .CLK(net116),
    .Q(\u_cpu.rf_ram.memory[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12348_ (.D(_01027_),
    .CLK(net117),
    .Q(\u_cpu.rf_ram.memory[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12349_ (.D(_01028_),
    .CLK(net125),
    .Q(\u_cpu.rf_ram.memory[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12350_ (.D(_01029_),
    .CLK(net135),
    .Q(\u_cpu.rf_ram.memory[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12351_ (.D(_01030_),
    .CLK(net138),
    .Q(\u_cpu.rf_ram.memory[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12352_ (.D(_01031_),
    .CLK(net135),
    .Q(\u_cpu.rf_ram.memory[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12353_ (.D(_01032_),
    .CLK(net112),
    .Q(\u_cpu.rf_ram.memory[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12354_ (.D(_01033_),
    .CLK(net117),
    .Q(\u_cpu.rf_ram.memory[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12355_ (.D(_01034_),
    .CLK(net116),
    .Q(\u_cpu.rf_ram.memory[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12356_ (.D(_01035_),
    .CLK(net117),
    .Q(\u_cpu.rf_ram.memory[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12357_ (.D(_01036_),
    .CLK(net125),
    .Q(\u_cpu.rf_ram.memory[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12358_ (.D(_01037_),
    .CLK(net127),
    .Q(\u_cpu.rf_ram.memory[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12359_ (.D(_01038_),
    .CLK(net138),
    .Q(\u_cpu.rf_ram.memory[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12360_ (.D(_01039_),
    .CLK(net135),
    .Q(\u_cpu.rf_ram.memory[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12361_ (.D(_01040_),
    .CLK(net211),
    .Q(\u_cpu.rf_ram.memory[93][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12362_ (.D(_01041_),
    .CLK(net211),
    .Q(\u_cpu.rf_ram.memory[93][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12363_ (.D(_01042_),
    .CLK(net211),
    .Q(\u_cpu.rf_ram.memory[93][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12364_ (.D(_01043_),
    .CLK(net210),
    .Q(\u_cpu.rf_ram.memory[93][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12365_ (.D(_01044_),
    .CLK(net210),
    .Q(\u_cpu.rf_ram.memory[93][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12366_ (.D(_01045_),
    .CLK(net210),
    .Q(\u_cpu.rf_ram.memory[93][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12367_ (.D(_01046_),
    .CLK(net210),
    .Q(\u_cpu.rf_ram.memory[93][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12368_ (.D(_01047_),
    .CLK(net210),
    .Q(\u_cpu.rf_ram.memory[93][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12369_ (.D(_01048_),
    .CLK(net351),
    .Q(\u_cpu.cpu.immdec.imm11_7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12370_ (.D(_01049_),
    .CLK(net359),
    .Q(\u_cpu.cpu.immdec.imm11_7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12371_ (.D(_01050_),
    .CLK(net343),
    .Q(\u_cpu.cpu.immdec.imm11_7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12372_ (.D(_01051_),
    .CLK(net343),
    .Q(\u_cpu.cpu.immdec.imm11_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12373_ (.D(_01052_),
    .CLK(net344),
    .Q(\u_cpu.cpu.immdec.imm11_7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12374_ (.D(_01053_),
    .CLK(net74),
    .Q(\u_cpu.rf_ram.memory[97][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12375_ (.D(_01054_),
    .CLK(net74),
    .Q(\u_cpu.rf_ram.memory[97][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12376_ (.D(_01055_),
    .CLK(net79),
    .Q(\u_cpu.rf_ram.memory[97][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12377_ (.D(_01056_),
    .CLK(net74),
    .Q(\u_cpu.rf_ram.memory[97][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12378_ (.D(_01057_),
    .CLK(net79),
    .Q(\u_cpu.rf_ram.memory[97][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12379_ (.D(_01058_),
    .CLK(net79),
    .Q(\u_cpu.rf_ram.memory[97][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12380_ (.D(_01059_),
    .CLK(net80),
    .Q(\u_cpu.rf_ram.memory[97][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12381_ (.D(_01060_),
    .CLK(net76),
    .Q(\u_cpu.rf_ram.memory[97][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12382_ (.D(_01061_),
    .CLK(net196),
    .Q(\u_cpu.rf_ram.memory[94][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12383_ (.D(_01062_),
    .CLK(net195),
    .Q(\u_cpu.rf_ram.memory[94][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12384_ (.D(_01063_),
    .CLK(net195),
    .Q(\u_cpu.rf_ram.memory[94][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12385_ (.D(_01064_),
    .CLK(net195),
    .Q(\u_cpu.rf_ram.memory[94][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12386_ (.D(_01065_),
    .CLK(net195),
    .Q(\u_cpu.rf_ram.memory[94][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12387_ (.D(_01066_),
    .CLK(net195),
    .Q(\u_cpu.rf_ram.memory[94][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12388_ (.D(_01067_),
    .CLK(net196),
    .Q(\u_cpu.rf_ram.memory[94][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12389_ (.D(_01068_),
    .CLK(net196),
    .Q(\u_cpu.rf_ram.memory[94][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12390_ (.D(_01069_),
    .CLK(net200),
    .Q(\u_cpu.rf_ram.memory[95][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12391_ (.D(_01070_),
    .CLK(net198),
    .Q(\u_cpu.rf_ram.memory[95][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12392_ (.D(_01071_),
    .CLK(net198),
    .Q(\u_cpu.rf_ram.memory[95][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12393_ (.D(_01072_),
    .CLK(net198),
    .Q(\u_cpu.rf_ram.memory[95][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12394_ (.D(_01073_),
    .CLK(net198),
    .Q(\u_cpu.rf_ram.memory[95][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12395_ (.D(_01074_),
    .CLK(net198),
    .Q(\u_cpu.rf_ram.memory[95][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12396_ (.D(_01075_),
    .CLK(net199),
    .Q(\u_cpu.rf_ram.memory[95][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12397_ (.D(_01076_),
    .CLK(net200),
    .Q(\u_cpu.rf_ram.memory[95][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12398_ (.D(_01077_),
    .CLK(net44),
    .Q(\u_cpu.rf_ram.memory[96][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12399_ (.D(_01078_),
    .CLK(net44),
    .Q(\u_cpu.rf_ram.memory[96][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12400_ (.D(_01079_),
    .CLK(net44),
    .Q(\u_cpu.rf_ram.memory[96][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12401_ (.D(_01080_),
    .CLK(net75),
    .Q(\u_cpu.rf_ram.memory[96][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12402_ (.D(_01081_),
    .CLK(net75),
    .Q(\u_cpu.rf_ram.memory[96][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12403_ (.D(_01082_),
    .CLK(net74),
    .Q(\u_cpu.rf_ram.memory[96][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12404_ (.D(_01083_),
    .CLK(net74),
    .Q(\u_cpu.rf_ram.memory[96][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12405_ (.D(_01084_),
    .CLK(net75),
    .Q(\u_cpu.rf_ram.memory[96][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12406_ (.D(_01085_),
    .CLK(net383),
    .Q(\u_cpu.cpu.bufreg.i_sh_signed ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12407_ (.D(_01086_),
    .CLK(net500),
    .Q(\u_cpu.cpu.genblk1.align.ctrl_misal ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12408_ (.D(_01087_),
    .CLK(net81),
    .Q(\u_cpu.rf_ram.memory[28][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12409_ (.D(_01088_),
    .CLK(net81),
    .Q(\u_cpu.rf_ram.memory[28][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12410_ (.D(_01089_),
    .CLK(net90),
    .Q(\u_cpu.rf_ram.memory[28][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12411_ (.D(_01090_),
    .CLK(net90),
    .Q(\u_cpu.rf_ram.memory[28][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12412_ (.D(_01091_),
    .CLK(net81),
    .Q(\u_cpu.rf_ram.memory[28][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12413_ (.D(_01092_),
    .CLK(net90),
    .Q(\u_cpu.rf_ram.memory[28][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12414_ (.D(_01093_),
    .CLK(net82),
    .Q(\u_cpu.rf_ram.memory[28][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12415_ (.D(_01094_),
    .CLK(net82),
    .Q(\u_cpu.rf_ram.memory[28][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12416_ (.D(_01095_),
    .CLK(net357),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12417_ (.D(_01096_),
    .CLK(net357),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12418_ (.D(_01097_),
    .CLK(net264),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12419_ (.D(_01098_),
    .CLK(net357),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12420_ (.D(_01099_),
    .CLK(net264),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12421_ (.D(_01100_),
    .CLK(net358),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12422_ (.D(_01101_),
    .CLK(net363),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12423_ (.D(_01102_),
    .CLK(net357),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12424_ (.D(_01103_),
    .CLK(net357),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12425_ (.D(_01104_),
    .CLK(net363),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12426_ (.D(_01105_),
    .CLK(net364),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12427_ (.D(_01106_),
    .CLK(net364),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12428_ (.D(_01107_),
    .CLK(net364),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12429_ (.D(_01108_),
    .CLK(net363),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12430_ (.D(_01109_),
    .CLK(net363),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12431_ (.D(_01110_),
    .CLK(net358),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12432_ (.D(_01111_),
    .CLK(net88),
    .Q(\u_cpu.rf_ram.memory[101][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12433_ (.D(_01112_),
    .CLK(net160),
    .Q(\u_cpu.rf_ram.memory[101][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12434_ (.D(_01113_),
    .CLK(net87),
    .Q(\u_cpu.rf_ram.memory[101][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12435_ (.D(_01114_),
    .CLK(net160),
    .Q(\u_cpu.rf_ram.memory[101][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12436_ (.D(_01115_),
    .CLK(net160),
    .Q(\u_cpu.rf_ram.memory[101][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12437_ (.D(_01116_),
    .CLK(net85),
    .Q(\u_cpu.rf_ram.memory[101][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12438_ (.D(_01117_),
    .CLK(net85),
    .Q(\u_cpu.rf_ram.memory[101][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12439_ (.D(_01118_),
    .CLK(net85),
    .Q(\u_cpu.rf_ram.memory[101][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12440_ (.D(_01119_),
    .CLK(net77),
    .Q(\u_cpu.rf_ram.memory[102][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12441_ (.D(_01120_),
    .CLK(net77),
    .Q(\u_cpu.rf_ram.memory[102][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12442_ (.D(_01121_),
    .CLK(net76),
    .Q(\u_cpu.rf_ram.memory[102][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12443_ (.D(_01122_),
    .CLK(net76),
    .Q(\u_cpu.rf_ram.memory[102][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12444_ (.D(_01123_),
    .CLK(net76),
    .Q(\u_cpu.rf_ram.memory[102][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12445_ (.D(_01124_),
    .CLK(net76),
    .Q(\u_cpu.rf_ram.memory[102][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12446_ (.D(_01125_),
    .CLK(net77),
    .Q(\u_cpu.rf_ram.memory[102][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12447_ (.D(_01126_),
    .CLK(net77),
    .Q(\u_cpu.rf_ram.memory[102][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12448_ (.D(_01127_),
    .CLK(net88),
    .Q(\u_cpu.rf_ram.memory[103][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12449_ (.D(_01128_),
    .CLK(net88),
    .Q(\u_cpu.rf_ram.memory[103][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12450_ (.D(_01129_),
    .CLK(net87),
    .Q(\u_cpu.rf_ram.memory[103][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12451_ (.D(_01130_),
    .CLK(net87),
    .Q(\u_cpu.rf_ram.memory[103][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12452_ (.D(_01131_),
    .CLK(net87),
    .Q(\u_cpu.rf_ram.memory[103][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12453_ (.D(_01132_),
    .CLK(net85),
    .Q(\u_cpu.rf_ram.memory[103][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12454_ (.D(_01133_),
    .CLK(net85),
    .Q(\u_cpu.rf_ram.memory[103][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12455_ (.D(_01134_),
    .CLK(net86),
    .Q(\u_cpu.rf_ram.memory[103][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12456_ (.D(_01135_),
    .CLK(net45),
    .Q(\u_cpu.rf_ram.memory[104][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12457_ (.D(_01136_),
    .CLK(net45),
    .Q(\u_cpu.rf_ram.memory[104][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12458_ (.D(_01137_),
    .CLK(net37),
    .Q(\u_cpu.rf_ram.memory[104][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12459_ (.D(_01138_),
    .CLK(net37),
    .Q(\u_cpu.rf_ram.memory[104][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12460_ (.D(_01139_),
    .CLK(net45),
    .Q(\u_cpu.rf_ram.memory[104][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12461_ (.D(_01140_),
    .CLK(net37),
    .Q(\u_cpu.rf_ram.memory[104][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12462_ (.D(_01141_),
    .CLK(net43),
    .Q(\u_cpu.rf_ram.memory[104][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12463_ (.D(_01142_),
    .CLK(net48),
    .Q(\u_cpu.rf_ram.memory[104][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12464_ (.D(_01143_),
    .CLK(net44),
    .Q(\u_cpu.rf_ram.memory[99][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12465_ (.D(_01144_),
    .CLK(net44),
    .Q(\u_cpu.rf_ram.memory[99][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12466_ (.D(_01145_),
    .CLK(net46),
    .Q(\u_cpu.rf_ram.memory[99][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12467_ (.D(_01146_),
    .CLK(net45),
    .Q(\u_cpu.rf_ram.memory[99][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12468_ (.D(_01147_),
    .CLK(net46),
    .Q(\u_cpu.rf_ram.memory[99][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12469_ (.D(_01148_),
    .CLK(net46),
    .Q(\u_cpu.rf_ram.memory[99][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12470_ (.D(_01149_),
    .CLK(net46),
    .Q(\u_cpu.rf_ram.memory[99][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12471_ (.D(_01150_),
    .CLK(net46),
    .Q(\u_cpu.rf_ram.memory[99][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12472_ (.D(_01151_),
    .CLK(net241),
    .Q(\u_cpu.rf_ram.memory[79][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12473_ (.D(_01152_),
    .CLK(net241),
    .Q(\u_cpu.rf_ram.memory[79][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12474_ (.D(_01153_),
    .CLK(net182),
    .Q(\u_cpu.rf_ram.memory[79][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12475_ (.D(_01154_),
    .CLK(net232),
    .Q(\u_cpu.rf_ram.memory[79][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12476_ (.D(_01155_),
    .CLK(net234),
    .Q(\u_cpu.rf_ram.memory[79][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12477_ (.D(_01156_),
    .CLK(net190),
    .Q(\u_cpu.rf_ram.memory[79][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12478_ (.D(_01157_),
    .CLK(net190),
    .Q(\u_cpu.rf_ram.memory[79][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12479_ (.D(_01158_),
    .CLK(net242),
    .Q(\u_cpu.rf_ram.memory[79][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12480_ (.D(_01159_),
    .CLK(net48),
    .Q(\u_cpu.rf_ram.memory[105][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12481_ (.D(_01160_),
    .CLK(net48),
    .Q(\u_cpu.rf_ram.memory[105][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12482_ (.D(_01161_),
    .CLK(net40),
    .Q(\u_cpu.rf_ram.memory[105][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12483_ (.D(_01162_),
    .CLK(net40),
    .Q(\u_cpu.rf_ram.memory[105][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12484_ (.D(_01163_),
    .CLK(net40),
    .Q(\u_cpu.rf_ram.memory[105][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12485_ (.D(_01164_),
    .CLK(net41),
    .Q(\u_cpu.rf_ram.memory[105][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12486_ (.D(_01165_),
    .CLK(net39),
    .Q(\u_cpu.rf_ram.memory[105][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12487_ (.D(_01166_),
    .CLK(net48),
    .Q(\u_cpu.rf_ram.memory[105][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12488_ (.D(_01167_),
    .CLK(net41),
    .Q(\u_cpu.rf_ram.memory[106][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12489_ (.D(_01168_),
    .CLK(net40),
    .Q(\u_cpu.rf_ram.memory[106][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12490_ (.D(_01169_),
    .CLK(net38),
    .Q(\u_cpu.rf_ram.memory[106][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12491_ (.D(_01170_),
    .CLK(net38),
    .Q(\u_cpu.rf_ram.memory[106][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12492_ (.D(_01171_),
    .CLK(net38),
    .Q(\u_cpu.rf_ram.memory[106][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12493_ (.D(_01172_),
    .CLK(net38),
    .Q(\u_cpu.rf_ram.memory[106][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12494_ (.D(_01173_),
    .CLK(net39),
    .Q(\u_cpu.rf_ram.memory[106][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12495_ (.D(_01174_),
    .CLK(net41),
    .Q(\u_cpu.rf_ram.memory[106][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12496_ (.D(_01175_),
    .CLK(net41),
    .Q(\u_cpu.rf_ram.memory[107][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12497_ (.D(_01176_),
    .CLK(net40),
    .Q(\u_cpu.rf_ram.memory[107][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12498_ (.D(_01177_),
    .CLK(net38),
    .Q(\u_cpu.rf_ram.memory[107][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12499_ (.D(_01178_),
    .CLK(net37),
    .Q(\u_cpu.rf_ram.memory[107][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12500_ (.D(_01179_),
    .CLK(net37),
    .Q(\u_cpu.rf_ram.memory[107][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12501_ (.D(_01180_),
    .CLK(net39),
    .Q(\u_cpu.rf_ram.memory[107][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12502_ (.D(_01181_),
    .CLK(net39),
    .Q(\u_cpu.rf_ram.memory[107][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12503_ (.D(_01182_),
    .CLK(net41),
    .Q(\u_cpu.rf_ram.memory[107][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12504_ (.D(_01183_),
    .CLK(net185),
    .Q(\u_cpu.rf_ram.memory[83][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12505_ (.D(_01184_),
    .CLK(net168),
    .Q(\u_cpu.rf_ram.memory[83][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12506_ (.D(_01185_),
    .CLK(net163),
    .Q(\u_cpu.rf_ram.memory[83][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12507_ (.D(_01186_),
    .CLK(net163),
    .Q(\u_cpu.rf_ram.memory[83][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12508_ (.D(_01187_),
    .CLK(net162),
    .Q(\u_cpu.rf_ram.memory[83][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12509_ (.D(_01188_),
    .CLK(net170),
    .Q(\u_cpu.rf_ram.memory[83][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12510_ (.D(_01189_),
    .CLK(net168),
    .Q(\u_cpu.rf_ram.memory[83][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12511_ (.D(_01190_),
    .CLK(net169),
    .Q(\u_cpu.rf_ram.memory[83][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12512_ (.D(_01191_),
    .CLK(net203),
    .Q(\u_cpu.rf_ram.memory[108][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12513_ (.D(_01192_),
    .CLK(net203),
    .Q(\u_cpu.rf_ram.memory[108][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12514_ (.D(_01193_),
    .CLK(net196),
    .Q(\u_cpu.rf_ram.memory[108][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12515_ (.D(_01194_),
    .CLK(net197),
    .Q(\u_cpu.rf_ram.memory[108][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12516_ (.D(_01195_),
    .CLK(net197),
    .Q(\u_cpu.rf_ram.memory[108][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12517_ (.D(_01196_),
    .CLK(net203),
    .Q(\u_cpu.rf_ram.memory[108][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12518_ (.D(_01197_),
    .CLK(net203),
    .Q(\u_cpu.rf_ram.memory[108][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12519_ (.D(_01198_),
    .CLK(net171),
    .Q(\u_cpu.rf_ram.memory[108][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12520_ (.D(_01199_),
    .CLK(net296),
    .Q(\u_cpu.rf_ram.memory[69][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12521_ (.D(_01200_),
    .CLK(net296),
    .Q(\u_cpu.rf_ram.memory[69][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12522_ (.D(_01201_),
    .CLK(net346),
    .Q(\u_cpu.rf_ram.memory[69][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12523_ (.D(_01202_),
    .CLK(net346),
    .Q(\u_cpu.rf_ram.memory[69][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12524_ (.D(_01203_),
    .CLK(net346),
    .Q(\u_cpu.rf_ram.memory[69][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12525_ (.D(_01204_),
    .CLK(net345),
    .Q(\u_cpu.rf_ram.memory[69][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12526_ (.D(_01205_),
    .CLK(net339),
    .Q(\u_cpu.rf_ram.memory[69][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12527_ (.D(_01206_),
    .CLK(net339),
    .Q(\u_cpu.rf_ram.memory[69][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12528_ (.D(_01207_),
    .CLK(net276),
    .Q(\u_cpu.rf_ram.memory[84][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12529_ (.D(_01208_),
    .CLK(net276),
    .Q(\u_cpu.rf_ram.memory[84][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12530_ (.D(_01209_),
    .CLK(net276),
    .Q(\u_cpu.rf_ram.memory[84][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12531_ (.D(_01210_),
    .CLK(net271),
    .Q(\u_cpu.rf_ram.memory[84][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12532_ (.D(_01211_),
    .CLK(net275),
    .Q(\u_cpu.rf_ram.memory[84][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12533_ (.D(_01212_),
    .CLK(net276),
    .Q(\u_cpu.rf_ram.memory[84][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12534_ (.D(_01213_),
    .CLK(net276),
    .Q(\u_cpu.rf_ram.memory[84][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12535_ (.D(_01214_),
    .CLK(net277),
    .Q(\u_cpu.rf_ram.memory[84][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12536_ (.D(_01215_),
    .CLK(net278),
    .Q(\u_cpu.rf_ram.memory[59][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12537_ (.D(_01216_),
    .CLK(net278),
    .Q(\u_cpu.rf_ram.memory[59][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12538_ (.D(_01217_),
    .CLK(net279),
    .Q(\u_cpu.rf_ram.memory[59][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12539_ (.D(_01218_),
    .CLK(net293),
    .Q(\u_cpu.rf_ram.memory[59][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12540_ (.D(_01219_),
    .CLK(net293),
    .Q(\u_cpu.rf_ram.memory[59][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12541_ (.D(_01220_),
    .CLK(net293),
    .Q(\u_cpu.rf_ram.memory[59][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12542_ (.D(_01221_),
    .CLK(net277),
    .Q(\u_cpu.rf_ram.memory[59][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12543_ (.D(_01222_),
    .CLK(net291),
    .Q(\u_cpu.rf_ram.memory[59][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12544_ (.D(_01223_),
    .CLK(net126),
    .Q(\u_cpu.rf_ram.memory[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12545_ (.D(_01224_),
    .CLK(net118),
    .Q(\u_cpu.rf_ram.memory[10][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12546_ (.D(_01225_),
    .CLK(net116),
    .Q(\u_cpu.rf_ram.memory[10][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12547_ (.D(_01226_),
    .CLK(net119),
    .Q(\u_cpu.rf_ram.memory[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12548_ (.D(_01227_),
    .CLK(net126),
    .Q(\u_cpu.rf_ram.memory[10][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12549_ (.D(_01228_),
    .CLK(net127),
    .Q(\u_cpu.rf_ram.memory[10][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12550_ (.D(_01229_),
    .CLK(net143),
    .Q(\u_cpu.rf_ram.memory[10][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12551_ (.D(_01230_),
    .CLK(net135),
    .Q(\u_cpu.rf_ram.memory[10][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12552_ (.D(_01231_),
    .CLK(net212),
    .Q(\u_cpu.rf_ram.memory[85][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12553_ (.D(_01232_),
    .CLK(net212),
    .Q(\u_cpu.rf_ram.memory[85][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12554_ (.D(_01233_),
    .CLK(net212),
    .Q(\u_cpu.rf_ram.memory[85][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12555_ (.D(_01234_),
    .CLK(net211),
    .Q(\u_cpu.rf_ram.memory[85][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12556_ (.D(_01235_),
    .CLK(net213),
    .Q(\u_cpu.rf_ram.memory[85][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12557_ (.D(_01236_),
    .CLK(net212),
    .Q(\u_cpu.rf_ram.memory[85][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12558_ (.D(_01237_),
    .CLK(net212),
    .Q(\u_cpu.rf_ram.memory[85][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12559_ (.D(_01238_),
    .CLK(net213),
    .Q(\u_cpu.rf_ram.memory[85][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12560_ (.D(_01239_),
    .CLK(net162),
    .Q(\u_cpu.rf_ram.memory[110][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12561_ (.D(_01240_),
    .CLK(net162),
    .Q(\u_cpu.rf_ram.memory[110][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12562_ (.D(_01241_),
    .CLK(net159),
    .Q(\u_cpu.rf_ram.memory[110][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12563_ (.D(_01242_),
    .CLK(net159),
    .Q(\u_cpu.rf_ram.memory[110][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12564_ (.D(_01243_),
    .CLK(net161),
    .Q(\u_cpu.rf_ram.memory[110][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12565_ (.D(_01244_),
    .CLK(net162),
    .Q(\u_cpu.rf_ram.memory[110][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12566_ (.D(_01245_),
    .CLK(net162),
    .Q(\u_cpu.rf_ram.memory[110][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12567_ (.D(_01246_),
    .CLK(net163),
    .Q(\u_cpu.rf_ram.memory[110][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12568_ (.D(_01247_),
    .CLK(net204),
    .Q(\u_cpu.rf_ram.memory[86][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12569_ (.D(_01248_),
    .CLK(net204),
    .Q(\u_cpu.rf_ram.memory[86][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12570_ (.D(_01249_),
    .CLK(net205),
    .Q(\u_cpu.rf_ram.memory[86][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12571_ (.D(_01250_),
    .CLK(net200),
    .Q(\u_cpu.rf_ram.memory[86][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12572_ (.D(_01251_),
    .CLK(net200),
    .Q(\u_cpu.rf_ram.memory[86][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12573_ (.D(_01252_),
    .CLK(net205),
    .Q(\u_cpu.rf_ram.memory[86][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12574_ (.D(_01253_),
    .CLK(net205),
    .Q(\u_cpu.rf_ram.memory[86][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12575_ (.D(_01254_),
    .CLK(net203),
    .Q(\u_cpu.rf_ram.memory[86][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12576_ (.D(_01255_),
    .CLK(net168),
    .Q(\u_cpu.rf_ram.memory[111][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12577_ (.D(_01256_),
    .CLK(net168),
    .Q(\u_cpu.rf_ram.memory[111][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12578_ (.D(_01257_),
    .CLK(net172),
    .Q(\u_cpu.rf_ram.memory[111][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12579_ (.D(_01258_),
    .CLK(net166),
    .Q(\u_cpu.rf_ram.memory[111][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12580_ (.D(_01259_),
    .CLK(net166),
    .Q(\u_cpu.rf_ram.memory[111][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12581_ (.D(_01260_),
    .CLK(net168),
    .Q(\u_cpu.rf_ram.memory[111][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12582_ (.D(_01261_),
    .CLK(net171),
    .Q(\u_cpu.rf_ram.memory[111][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12583_ (.D(_01262_),
    .CLK(net169),
    .Q(\u_cpu.rf_ram.memory[111][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12584_ (.D(_01263_),
    .CLK(net207),
    .Q(\u_cpu.rf_ram.memory[87][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12585_ (.D(_01264_),
    .CLK(net207),
    .Q(\u_cpu.rf_ram.memory[87][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12586_ (.D(_01265_),
    .CLK(net205),
    .Q(\u_cpu.rf_ram.memory[87][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12587_ (.D(_01266_),
    .CLK(net200),
    .Q(\u_cpu.rf_ram.memory[87][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12588_ (.D(_01267_),
    .CLK(net201),
    .Q(\u_cpu.rf_ram.memory[87][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12589_ (.D(_01268_),
    .CLK(net205),
    .Q(\u_cpu.rf_ram.memory[87][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12590_ (.D(_01269_),
    .CLK(net206),
    .Q(\u_cpu.rf_ram.memory[87][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12591_ (.D(_01270_),
    .CLK(net206),
    .Q(\u_cpu.rf_ram.memory[87][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12592_ (.D(_01271_),
    .CLK(net278),
    .Q(\u_cpu.rf_ram.memory[88][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12593_ (.D(_01272_),
    .CLK(net278),
    .Q(\u_cpu.rf_ram.memory[88][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12594_ (.D(_01273_),
    .CLK(net279),
    .Q(\u_cpu.rf_ram.memory[88][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12595_ (.D(_01274_),
    .CLK(net274),
    .Q(\u_cpu.rf_ram.memory[88][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12596_ (.D(_01275_),
    .CLK(net274),
    .Q(\u_cpu.rf_ram.memory[88][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12597_ (.D(_01276_),
    .CLK(net279),
    .Q(\u_cpu.rf_ram.memory[88][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12598_ (.D(_01277_),
    .CLK(net279),
    .Q(\u_cpu.rf_ram.memory[88][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12599_ (.D(_01278_),
    .CLK(net278),
    .Q(\u_cpu.rf_ram.memory[88][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12600_ (.D(_01279_),
    .CLK(net378),
    .Q(\u_cpu.cpu.genblk3.csr.mcause3_0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12601_ (.D(_01280_),
    .CLK(net374),
    .Q(\u_cpu.cpu.genblk3.csr.mcause3_0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12602_ (.D(_01281_),
    .CLK(net373),
    .Q(\u_cpu.cpu.genblk3.csr.mcause3_0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12603_ (.D(_01282_),
    .CLK(net374),
    .Q(\u_cpu.cpu.genblk3.csr.mcause3_0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12604_ (.D(_01283_),
    .CLK(net378),
    .Q(\u_cpu.cpu.genblk3.csr.mcause31 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12605_ (.D(_01284_),
    .CLK(net378),
    .Q(\u_cpu.cpu.genblk3.csr.mstatus_mpie ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12606_ (.D(_01285_),
    .CLK(net480),
    .Q(\u_cpu.cpu.genblk3.csr.mie_mtie ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12607_ (.D(_01286_),
    .CLK(net380),
    .Q(\u_cpu.cpu.genblk3.csr.mstatus_mie ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12608_ (.D(_01287_),
    .CLK(net360),
    .Q(\u_cpu.cpu.ctrl.i_iscomp ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12609_ (.D(_01288_),
    .CLK(net380),
    .Q(\u_cpu.cpu.genblk3.csr.o_new_irq ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12610_ (.D(_01289_),
    .CLK(net52),
    .Q(\u_cpu.rf_ram.memory[27][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12611_ (.D(_01290_),
    .CLK(net52),
    .Q(\u_cpu.rf_ram.memory[27][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12612_ (.D(_01291_),
    .CLK(net51),
    .Q(\u_cpu.rf_ram.memory[27][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12613_ (.D(_01292_),
    .CLK(net51),
    .Q(\u_cpu.rf_ram.memory[27][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12614_ (.D(_01293_),
    .CLK(net51),
    .Q(\u_cpu.rf_ram.memory[27][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12615_ (.D(_01294_),
    .CLK(net56),
    .Q(\u_cpu.rf_ram.memory[27][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12616_ (.D(_01295_),
    .CLK(net56),
    .Q(\u_cpu.rf_ram.memory[27][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12617_ (.D(_01296_),
    .CLK(net56),
    .Q(\u_cpu.rf_ram.memory[27][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12618_ (.D(_01297_),
    .CLK(net52),
    .Q(\u_cpu.rf_ram.memory[26][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12619_ (.D(_01298_),
    .CLK(net52),
    .Q(\u_cpu.rf_ram.memory[26][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12620_ (.D(_01299_),
    .CLK(net51),
    .Q(\u_cpu.rf_ram.memory[26][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12621_ (.D(_01300_),
    .CLK(net51),
    .Q(\u_cpu.rf_ram.memory[26][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12622_ (.D(_01301_),
    .CLK(net53),
    .Q(\u_cpu.rf_ram.memory[26][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12623_ (.D(_01302_),
    .CLK(net52),
    .Q(\u_cpu.rf_ram.memory[26][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12624_ (.D(_01303_),
    .CLK(net57),
    .Q(\u_cpu.rf_ram.memory[26][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12625_ (.D(_01304_),
    .CLK(net57),
    .Q(\u_cpu.rf_ram.memory[26][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12626_ (.D(_01305_),
    .CLK(net53),
    .Q(\u_cpu.rf_ram.memory[25][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12627_ (.D(_01306_),
    .CLK(net54),
    .Q(\u_cpu.rf_ram.memory[25][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12628_ (.D(_01307_),
    .CLK(net53),
    .Q(\u_cpu.rf_ram.memory[25][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12629_ (.D(_01308_),
    .CLK(net53),
    .Q(\u_cpu.rf_ram.memory[25][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12630_ (.D(_01309_),
    .CLK(net53),
    .Q(\u_cpu.rf_ram.memory[25][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12631_ (.D(_01310_),
    .CLK(net59),
    .Q(\u_cpu.rf_ram.memory[25][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12632_ (.D(_01311_),
    .CLK(net59),
    .Q(\u_cpu.rf_ram.memory[25][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12633_ (.D(_01312_),
    .CLK(net54),
    .Q(\u_cpu.rf_ram.memory[25][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12634_ (.D(_01313_),
    .CLK(net63),
    .Q(\u_cpu.rf_ram.memory[24][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12635_ (.D(_01314_),
    .CLK(net63),
    .Q(\u_cpu.rf_ram.memory[24][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12636_ (.D(_01315_),
    .CLK(net63),
    .Q(\u_cpu.rf_ram.memory[24][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12637_ (.D(_01316_),
    .CLK(net63),
    .Q(\u_cpu.rf_ram.memory[24][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12638_ (.D(_01317_),
    .CLK(net63),
    .Q(\u_cpu.rf_ram.memory[24][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12639_ (.D(_01318_),
    .CLK(net64),
    .Q(\u_cpu.rf_ram.memory[24][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12640_ (.D(_01319_),
    .CLK(net67),
    .Q(\u_cpu.rf_ram.memory[24][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12641_ (.D(_01320_),
    .CLK(net64),
    .Q(\u_cpu.rf_ram.memory[24][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12642_ (.D(_01321_),
    .CLK(net112),
    .Q(\u_cpu.rf_ram.memory[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12643_ (.D(_01322_),
    .CLK(net115),
    .Q(\u_cpu.rf_ram.memory[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12644_ (.D(_01323_),
    .CLK(net113),
    .Q(\u_cpu.rf_ram.memory[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12645_ (.D(_01324_),
    .CLK(net124),
    .Q(\u_cpu.rf_ram.memory[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12646_ (.D(_01325_),
    .CLK(net123),
    .Q(\u_cpu.rf_ram.memory[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12647_ (.D(_01326_),
    .CLK(net133),
    .Q(\u_cpu.rf_ram.memory[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12648_ (.D(_01327_),
    .CLK(net142),
    .Q(\u_cpu.rf_ram.memory[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12649_ (.D(_01328_),
    .CLK(net134),
    .Q(\u_cpu.rf_ram.memory[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12650_ (.D(_01329_),
    .CLK(net65),
    .Q(\u_cpu.rf_ram.memory[98][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12651_ (.D(_01330_),
    .CLK(net65),
    .Q(\u_cpu.rf_ram.memory[98][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12652_ (.D(_01331_),
    .CLK(net66),
    .Q(\u_cpu.rf_ram.memory[98][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12653_ (.D(_01332_),
    .CLK(net66),
    .Q(\u_cpu.rf_ram.memory[98][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12654_ (.D(_01333_),
    .CLK(net93),
    .Q(\u_cpu.rf_ram.memory[98][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12655_ (.D(_01334_),
    .CLK(net47),
    .Q(\u_cpu.rf_ram.memory[98][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12656_ (.D(_01335_),
    .CLK(net47),
    .Q(\u_cpu.rf_ram.memory[98][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12657_ (.D(_01336_),
    .CLK(net80),
    .Q(\u_cpu.rf_ram.memory[98][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12658_ (.D(_01337_),
    .CLK(net160),
    .Q(\u_cpu.rf_ram.memory[100][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12659_ (.D(_01338_),
    .CLK(net160),
    .Q(\u_cpu.rf_ram.memory[100][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12660_ (.D(_01339_),
    .CLK(net159),
    .Q(\u_cpu.rf_ram.memory[100][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12661_ (.D(_01340_),
    .CLK(net159),
    .Q(\u_cpu.rf_ram.memory[100][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12662_ (.D(_01341_),
    .CLK(net159),
    .Q(\u_cpu.rf_ram.memory[100][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12663_ (.D(_01342_),
    .CLK(net87),
    .Q(\u_cpu.rf_ram.memory[100][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12664_ (.D(_01343_),
    .CLK(net86),
    .Q(\u_cpu.rf_ram.memory[100][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12665_ (.D(_01344_),
    .CLK(net88),
    .Q(\u_cpu.rf_ram.memory[100][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12666_ (.D(_01345_),
    .CLK(net286),
    .Q(\u_cpu.rf_ram.memory[89][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12667_ (.D(_01346_),
    .CLK(net287),
    .Q(\u_cpu.rf_ram.memory[89][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12668_ (.D(_01347_),
    .CLK(net286),
    .Q(\u_cpu.rf_ram.memory[89][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12669_ (.D(_01348_),
    .CLK(net286),
    .Q(\u_cpu.rf_ram.memory[89][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12670_ (.D(_01349_),
    .CLK(net286),
    .Q(\u_cpu.rf_ram.memory[89][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12671_ (.D(_01350_),
    .CLK(net288),
    .Q(\u_cpu.rf_ram.memory[89][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12672_ (.D(_01351_),
    .CLK(net288),
    .Q(\u_cpu.rf_ram.memory[89][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12673_ (.D(_01352_),
    .CLK(net289),
    .Q(\u_cpu.rf_ram.memory[89][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12674_ (.D(_00025_),
    .CLK(net256),
    .Q(\u_cpu.rf_ram.regzero ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12675_ (.D(_01353_),
    .CLK(net102),
    .Q(\u_cpu.rf_ram.memory[23][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12676_ (.D(_01354_),
    .CLK(net102),
    .Q(\u_cpu.rf_ram.memory[23][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12677_ (.D(_01355_),
    .CLK(net95),
    .Q(\u_cpu.rf_ram.memory[23][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12678_ (.D(_01356_),
    .CLK(net95),
    .Q(\u_cpu.rf_ram.memory[23][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12679_ (.D(_01357_),
    .CLK(net96),
    .Q(\u_cpu.rf_ram.memory[23][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12680_ (.D(_01358_),
    .CLK(net96),
    .Q(\u_cpu.rf_ram.memory[23][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12681_ (.D(_01359_),
    .CLK(net97),
    .Q(\u_cpu.rf_ram.memory[23][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12682_ (.D(_01360_),
    .CLK(net100),
    .Q(\u_cpu.rf_ram.memory[23][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12683_ (.D(_01361_),
    .CLK(net496),
    .Q(\u_cpu.cpu.state.ibus_cyc ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12684_ (.D(\u_cpu.rf_ram_if.wdata0_r[1] ),
    .CLK(net232),
    .Q(\u_cpu.rf_ram_if.wdata0_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12685_ (.D(\u_cpu.rf_ram_if.wdata0_r[2] ),
    .CLK(net140),
    .Q(\u_cpu.rf_ram_if.wdata0_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12686_ (.D(\u_cpu.rf_ram_if.wdata0_r[3] ),
    .CLK(net232),
    .Q(\u_cpu.rf_ram_if.wdata0_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12687_ (.D(\u_cpu.rf_ram_if.wdata0_r[4] ),
    .CLK(net232),
    .Q(\u_cpu.rf_ram_if.wdata0_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12688_ (.D(\u_cpu.rf_ram_if.wdata0_r[5] ),
    .CLK(net234),
    .Q(\u_cpu.rf_ram_if.wdata0_r[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12689_ (.D(\u_cpu.rf_ram_if.wdata0_r[6] ),
    .CLK(net234),
    .Q(\u_cpu.rf_ram_if.wdata0_r[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12690_ (.D(\u_cpu.cpu.o_wdata0 ),
    .CLK(net234),
    .Q(\u_cpu.rf_ram_if.wdata0_r[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12691_ (.D(\u_cpu.rf_ram_if.wtrig0 ),
    .CLK(net342),
    .Q(\u_cpu.rf_ram_if.genblk1.wtrig0_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12692_ (.D(_01362_),
    .CLK(net252),
    .Q(\u_cpu.rf_ram_if.rdata1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12693_ (.D(_01363_),
    .CLK(net257),
    .Q(\u_cpu.rf_ram_if.rdata0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12694_ (.D(_01364_),
    .CLK(net379),
    .Q(\u_cpu.rf_ram_if.rgnt ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12695_ (.D(\u_cpu.rf_ram_if.rtrig0 ),
    .CLK(net260),
    .Q(\u_cpu.rf_ram_if.rtrig1 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12696_ (.D(_01365_),
    .CLK(net379),
    .Q(\u_cpu.rf_ram_if.rcnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12697_ (.D(\u_cpu.rf_ram_if.wdata1_r[1] ),
    .CLK(net140),
    .Q(\u_cpu.rf_ram_if.wdata1_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12698_ (.D(\u_cpu.rf_ram_if.wdata1_r[2] ),
    .CLK(net140),
    .Q(\u_cpu.rf_ram_if.wdata1_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12699_ (.D(\u_cpu.rf_ram_if.wdata1_r[3] ),
    .CLK(net232),
    .Q(\u_cpu.rf_ram_if.wdata1_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12700_ (.D(\u_cpu.rf_ram_if.wdata1_r[4] ),
    .CLK(net141),
    .Q(\u_cpu.rf_ram_if.wdata1_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12701_ (.D(\u_cpu.rf_ram_if.wdata1_r[5] ),
    .CLK(net233),
    .Q(\u_cpu.rf_ram_if.wdata1_r[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12702_ (.D(\u_cpu.rf_ram_if.wdata1_r[6] ),
    .CLK(net233),
    .Q(\u_cpu.rf_ram_if.wdata1_r[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12703_ (.D(\u_cpu.rf_ram_if.wdata1_r[7] ),
    .CLK(net235),
    .Q(\u_cpu.rf_ram_if.wdata1_r[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12704_ (.D(\u_cpu.cpu.o_wdata1 ),
    .CLK(net239),
    .Q(\u_cpu.rf_ram_if.wdata1_r[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12705_ (.D(\u_cpu.cpu.o_wen0 ),
    .CLK(net353),
    .Q(\u_cpu.rf_ram_if.wen0_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12706_ (.D(\u_cpu.cpu.o_wen1 ),
    .CLK(net353),
    .Q(\u_cpu.rf_ram_if.wen1_r ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06969__A1 (.I(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07121__A1 (.I(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11098__A2 (.I(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11116__B (.I(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05743__A3 (.I(_01393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11089__A2 (.I(_01393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11102__A2 (.I(_01393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05741__A1 (.I(_01391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06946__A2 (.I(_01391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10071__A1 (.I(_01391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05739__A2 (.I(_01389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05752__A2 (.I(_01389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05770__A2 (.I(_01389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05774__A2 (.I(_01389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05738__A3 (.I(_01388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05745__B (.I(_01388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05754__A2 (.I(_01388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05765__A2 (.I(_01388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07113__A1 (.I(_01388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05737__B (.I(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06970__I (.I(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07126__A1 (.I(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07127__A2 (.I(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05736__C (.I(_01386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06985__A3 (.I(_01386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07713__A2 (.I(_01386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11090__A1 (.I(_01386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11094__B2 (.I(_01386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05736__B (.I(_01385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06985__A1 (.I(_01385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05732__B (.I(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07029__B1 (.I(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09841__A1 (.I(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11102__A1 (.I(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05738__A2 (.I(_01378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05754__A1 (.I(_01378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05764__C (.I(_01378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11116__A2 (.I(_01378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05727__A3 (.I(_01377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05762__A2 (.I(_01377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09922__A3 (.I(_01377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05724__I (.I(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06988__B (.I(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07018__A1 (.I(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07083__I (.I(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07701__A1 (.I(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05722__A3 (.I(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05733__A4 (.I(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06949__I (.I(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06976__A1 (.I(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07122__A2 (.I(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05722__A2 (.I(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06948__I (.I(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06951__I (.I(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06987__A2 (.I(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06991__A2 (.I(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05715__I (.I(_01367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05745__C (.I(_01367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05750__I (.I(_01367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05769__A2 (.I(_01367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05773__A2 (.I(_01367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12371__D (.I(_01050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12205__D (.I(_00888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07016__A3 (.I(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12045__D (.I(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12674__D (.I(_00025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11750__D (.I(_00007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11749__D (.I(_00006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11748__D (.I(_00005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11747__D (.I(_00004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11746__D (.I(_00003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11745__D (.I(_00002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11744__D (.I(_00001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11743__D (.I(_00000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06527__A1 (.I(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05772__I (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06030__I (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06246__I (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06778__A1 (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06866__A1 (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05778__A2 (.I(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06217__B (.I(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06335__B (.I(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06448__B (.I(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06562__B (.I(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05768__I (.I(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06027__I (.I(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06153__I (.I(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06188__I (.I(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06455__I (.I(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05767__I (.I(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05970__I (.I(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06061__I (.I(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06106__I (.I(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06493__I (.I(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05764__A2 (.I(_01414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07132__A2 (.I(_01414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05764__A1 (.I(_01413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06958__A2 (.I(_01413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06964__A3 (.I(_01413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05762__A1 (.I(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06983__A1 (.I(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10358__A2 (.I(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05761__A2 (.I(_01411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06968__A1 (.I(_01411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06988__A1 (.I(_01411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07011__B2 (.I(_01411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07081__B1 (.I(_01411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05761__A1 (.I(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07710__A1 (.I(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09204__A1 (.I(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09825__A1 (.I(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05758__I (.I(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06945__I (.I(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06975__B (.I(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06987__A1 (.I(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06992__A2 (.I(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05778__A1 (.I(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05947__I (.I(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06741__A1 (.I(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06829__A1 (.I(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06917__A1 (.I(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05755__A2 (.I(_01405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06218__I (.I(_01405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06739__C (.I(_01405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06827__C (.I(_01405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06915__C (.I(_01405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05755__A1 (.I(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06193__I (.I(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06730__B (.I(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06818__B (.I(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06906__B (.I(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05751__A2 (.I(_01401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05754__B (.I(_01401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05780__I (.I(_01401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07063__I (.I(_01401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07068__I (.I(_01401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05779__A1 (.I(_01400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06201__A1 (.I(_01400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06328__A1 (.I(_01400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06440__A1 (.I(_01400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06554__A1 (.I(_01400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05747__I (.I(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05992__I (.I(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06031__I (.I(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06048__I (.I(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06160__I (.I(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__tiel serv_1_566 (.ZN(net566));
 gf180mcu_fd_sc_mcu7t5v0__tiel serv_1_567 (.ZN(net567));
 gf180mcu_fd_sc_mcu7t5v0__tiel serv_1_568 (.ZN(net568));
 gf180mcu_fd_sc_mcu7t5v0__tiel serv_1_569 (.ZN(net569));
 gf180mcu_fd_sc_mcu7t5v0__tiel serv_1_570 (.ZN(net570));
 gf180mcu_fd_sc_mcu7t5v0__tiel serv_1_571 (.ZN(net571));
 gf180mcu_fd_sc_mcu7t5v0__tiel serv_1_572 (.ZN(net572));
 gf180mcu_fd_sc_mcu7t5v0__tiel serv_1_573 (.ZN(net573));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05745__A1 (.I(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12863_ (.I(\u_scanchain_local.clk_out ),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12864_ (.I(\u_scanchain_local.data_out ),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \u_scanchain_local.input_buf_clk  (.I(net1),
    .Z(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__dffnq_1 \u_scanchain_local.out_flop  (.D(\u_scanchain_local.module_data_in[69] ),
    .CLKN(net26),
    .Q(\u_scanchain_local.data_out_i ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \u_scanchain_local.output_buffers[2]  (.I(\u_scanchain_local.data_out_i ),
    .Z(\u_scanchain_local.data_out ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \u_scanchain_local.output_buffers[3]  (.I(net34),
    .Z(\u_scanchain_local.clk_out ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[0]  (.D(net3),
    .SE(net552),
    .SI(\u_arbiter.o_wb_cpu_cyc ),
    .CLK(net20),
    .Q(\u_cpu.cpu.genblk3.csr.i_mtip ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[10]  (.D(\u_arbiter.i_wb_cpu_rdt[7] ),
    .SE(net544),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[4] ),
    .CLK(net12),
    .Q(\u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[11]  (.D(\u_arbiter.i_wb_cpu_rdt[8] ),
    .SE(net544),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .CLK(net12),
    .Q(\u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[12]  (.D(\u_arbiter.i_wb_cpu_rdt[9] ),
    .SE(net544),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[6] ),
    .CLK(net12),
    .Q(\u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[13]  (.D(\u_arbiter.i_wb_cpu_rdt[10] ),
    .SE(net544),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[7] ),
    .CLK(net12),
    .Q(\u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[14]  (.D(\u_arbiter.i_wb_cpu_rdt[11] ),
    .SE(net542),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[8] ),
    .CLK(net11),
    .Q(\u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[15]  (.D(\u_arbiter.i_wb_cpu_rdt[12] ),
    .SE(net542),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[9] ),
    .CLK(net11),
    .Q(\u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[16]  (.D(\u_arbiter.i_wb_cpu_rdt[13] ),
    .SE(net542),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[10] ),
    .CLK(net11),
    .Q(\u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[17]  (.D(\u_arbiter.i_wb_cpu_rdt[14] ),
    .SE(net542),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[11] ),
    .CLK(net11),
    .Q(\u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[18]  (.D(\u_arbiter.i_wb_cpu_rdt[15] ),
    .SE(net542),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[12] ),
    .CLK(net9),
    .Q(\u_arbiter.i_wb_cpu_rdt[16] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[19]  (.D(\u_arbiter.i_wb_cpu_rdt[16] ),
    .SE(net541),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[13] ),
    .CLK(net9),
    .Q(\u_arbiter.i_wb_cpu_rdt[17] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[1]  (.D(\u_cpu.cpu.genblk3.csr.i_mtip ),
    .SE(net552),
    .SI(\u_arbiter.o_wb_cpu_we ),
    .CLK(net20),
    .Q(\u_arbiter.i_wb_cpu_ack ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[20]  (.D(\u_arbiter.i_wb_cpu_rdt[17] ),
    .SE(net541),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[14] ),
    .CLK(net9),
    .Q(\u_arbiter.i_wb_cpu_rdt[18] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[21]  (.D(\u_arbiter.i_wb_cpu_rdt[18] ),
    .SE(net541),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[15] ),
    .CLK(net9),
    .Q(\u_arbiter.i_wb_cpu_rdt[19] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[22]  (.D(\u_arbiter.i_wb_cpu_rdt[19] ),
    .SE(net545),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[16] ),
    .CLK(net13),
    .Q(\u_arbiter.i_wb_cpu_rdt[20] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[23]  (.D(\u_arbiter.i_wb_cpu_rdt[20] ),
    .SE(net541),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[17] ),
    .CLK(net10),
    .Q(\u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[24]  (.D(\u_arbiter.i_wb_cpu_rdt[21] ),
    .SE(net541),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[18] ),
    .CLK(net9),
    .Q(\u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[25]  (.D(\u_arbiter.i_wb_cpu_rdt[22] ),
    .SE(net543),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[19] ),
    .CLK(net10),
    .Q(\u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[26]  (.D(\u_arbiter.i_wb_cpu_rdt[23] ),
    .SE(net545),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[20] ),
    .CLK(net13),
    .Q(\u_arbiter.i_wb_cpu_rdt[24] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[27]  (.D(\u_arbiter.i_wb_cpu_rdt[24] ),
    .SE(net547),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[21] ),
    .CLK(net13),
    .Q(\u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[28]  (.D(\u_arbiter.i_wb_cpu_rdt[25] ),
    .SE(net547),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[22] ),
    .CLK(net17),
    .Q(\u_arbiter.i_wb_cpu_rdt[26] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[29]  (.D(\u_arbiter.i_wb_cpu_rdt[26] ),
    .SE(net545),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[23] ),
    .CLK(net13),
    .Q(\u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[2]  (.D(net8),
    .SE(net548),
    .SI(\u_arbiter.i_wb_cpu_dbus_sel[0] ),
    .CLK(net15),
    .Q(\u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[30]  (.D(\u_arbiter.i_wb_cpu_rdt[27] ),
    .SE(net547),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[24] ),
    .CLK(net17),
    .Q(\u_arbiter.i_wb_cpu_rdt[28] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[31]  (.D(\u_arbiter.i_wb_cpu_rdt[28] ),
    .SE(net547),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[25] ),
    .CLK(net17),
    .Q(\u_arbiter.i_wb_cpu_rdt[29] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[32]  (.D(\u_arbiter.i_wb_cpu_rdt[29] ),
    .SE(net549),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[26] ),
    .CLK(net16),
    .Q(\u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[33]  (.D(\u_arbiter.i_wb_cpu_rdt[30] ),
    .SE(net550),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[27] ),
    .CLK(net17),
    .Q(\u_arbiter.i_wb_cpu_rdt[31] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[34]  (.D(\u_arbiter.i_wb_cpu_rdt[31] ),
    .SE(net549),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[28] ),
    .CLK(net16),
    .Q(\u_scanchain_local.module_data_in[34] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[35]  (.D(\u_scanchain_local.module_data_in[34] ),
    .SE(net549),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[29] ),
    .CLK(net16),
    .Q(\u_scanchain_local.module_data_in[35] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[36]  (.D(\u_scanchain_local.module_data_in[35] ),
    .SE(net556),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[30] ),
    .CLK(net24),
    .Q(\u_scanchain_local.module_data_in[36] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[37]  (.D(\u_scanchain_local.module_data_in[36] ),
    .SE(net556),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[31] ),
    .CLK(net24),
    .Q(\u_scanchain_local.module_data_in[37] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[38]  (.D(\u_scanchain_local.module_data_in[37] ),
    .SE(net552),
    .SI(\u_arbiter.o_wb_cpu_adr[0] ),
    .CLK(net20),
    .Q(\u_scanchain_local.module_data_in[38] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[39]  (.D(\u_scanchain_local.module_data_in[38] ),
    .SE(net552),
    .SI(\u_arbiter.o_wb_cpu_adr[1] ),
    .CLK(net20),
    .Q(\u_scanchain_local.module_data_in[39] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[3]  (.D(\u_arbiter.i_wb_cpu_rdt[0] ),
    .SE(net547),
    .SI(\u_arbiter.i_wb_cpu_dbus_sel[1] ),
    .CLK(net17),
    .Q(\u_arbiter.i_wb_cpu_rdt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[40]  (.D(\u_scanchain_local.module_data_in[39] ),
    .SE(net552),
    .SI(\u_arbiter.o_wb_cpu_adr[2] ),
    .CLK(net20),
    .Q(\u_scanchain_local.module_data_in[40] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[41]  (.D(\u_scanchain_local.module_data_in[40] ),
    .SE(net553),
    .SI(\u_arbiter.o_wb_cpu_adr[3] ),
    .CLK(net21),
    .Q(\u_scanchain_local.module_data_in[41] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[42]  (.D(\u_scanchain_local.module_data_in[41] ),
    .SE(net553),
    .SI(\u_arbiter.o_wb_cpu_adr[4] ),
    .CLK(net21),
    .Q(\u_scanchain_local.module_data_in[42] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[43]  (.D(\u_scanchain_local.module_data_in[42] ),
    .SE(net559),
    .SI(\u_arbiter.o_wb_cpu_adr[5] ),
    .CLK(net27),
    .Q(\u_scanchain_local.module_data_in[43] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[44]  (.D(\u_scanchain_local.module_data_in[43] ),
    .SE(net559),
    .SI(\u_arbiter.o_wb_cpu_adr[6] ),
    .CLK(net27),
    .Q(\u_scanchain_local.module_data_in[44] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[45]  (.D(\u_scanchain_local.module_data_in[44] ),
    .SE(net559),
    .SI(\u_arbiter.o_wb_cpu_adr[7] ),
    .CLK(net27),
    .Q(\u_scanchain_local.module_data_in[45] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[46]  (.D(\u_scanchain_local.module_data_in[45] ),
    .SE(net558),
    .SI(\u_arbiter.o_wb_cpu_adr[8] ),
    .CLK(net26),
    .Q(\u_scanchain_local.module_data_in[46] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[47]  (.D(\u_scanchain_local.module_data_in[46] ),
    .SE(net558),
    .SI(\u_arbiter.o_wb_cpu_adr[9] ),
    .CLK(net26),
    .Q(\u_scanchain_local.module_data_in[47] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[48]  (.D(\u_scanchain_local.module_data_in[47] ),
    .SE(net558),
    .SI(\u_arbiter.o_wb_cpu_adr[10] ),
    .CLK(net26),
    .Q(\u_scanchain_local.module_data_in[48] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[49]  (.D(\u_scanchain_local.module_data_in[48] ),
    .SE(net558),
    .SI(\u_arbiter.o_wb_cpu_adr[11] ),
    .CLK(net28),
    .Q(\u_scanchain_local.module_data_in[49] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[4]  (.D(\u_arbiter.i_wb_cpu_rdt[1] ),
    .SE(net548),
    .SI(\u_arbiter.i_wb_cpu_dbus_sel[2] ),
    .CLK(net15),
    .Q(\u_arbiter.i_wb_cpu_rdt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[50]  (.D(\u_scanchain_local.module_data_in[49] ),
    .SE(net558),
    .SI(\u_arbiter.o_wb_cpu_adr[12] ),
    .CLK(net26),
    .Q(\u_scanchain_local.module_data_in[50] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[51]  (.D(\u_scanchain_local.module_data_in[50] ),
    .SE(net560),
    .SI(\u_arbiter.o_wb_cpu_adr[13] ),
    .CLK(net29),
    .Q(\u_scanchain_local.module_data_in[51] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[52]  (.D(\u_scanchain_local.module_data_in[51] ),
    .SE(net561),
    .SI(\u_arbiter.o_wb_cpu_adr[14] ),
    .CLK(net29),
    .Q(\u_scanchain_local.module_data_in[52] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[53]  (.D(\u_scanchain_local.module_data_in[52] ),
    .SE(net561),
    .SI(\u_arbiter.o_wb_cpu_adr[15] ),
    .CLK(net29),
    .Q(\u_scanchain_local.module_data_in[53] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[54]  (.D(\u_scanchain_local.module_data_in[53] ),
    .SE(net561),
    .SI(\u_arbiter.o_wb_cpu_adr[16] ),
    .CLK(net29),
    .Q(\u_scanchain_local.module_data_in[54] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[55]  (.D(\u_scanchain_local.module_data_in[54] ),
    .SE(net561),
    .SI(\u_arbiter.o_wb_cpu_adr[17] ),
    .CLK(net29),
    .Q(\u_scanchain_local.module_data_in[55] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[56]  (.D(\u_scanchain_local.module_data_in[55] ),
    .SE(net561),
    .SI(\u_arbiter.o_wb_cpu_adr[18] ),
    .CLK(net30),
    .Q(\u_scanchain_local.module_data_in[56] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[57]  (.D(\u_scanchain_local.module_data_in[56] ),
    .SE(net562),
    .SI(\u_arbiter.o_wb_cpu_adr[19] ),
    .CLK(net31),
    .Q(\u_scanchain_local.module_data_in[57] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[58]  (.D(\u_scanchain_local.module_data_in[57] ),
    .SE(net562),
    .SI(\u_arbiter.o_wb_cpu_adr[20] ),
    .CLK(net30),
    .Q(\u_scanchain_local.module_data_in[58] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[59]  (.D(\u_scanchain_local.module_data_in[58] ),
    .SE(net562),
    .SI(\u_arbiter.o_wb_cpu_adr[21] ),
    .CLK(net31),
    .Q(\u_scanchain_local.module_data_in[59] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[5]  (.D(\u_arbiter.i_wb_cpu_rdt[2] ),
    .SE(net548),
    .SI(\u_arbiter.i_wb_cpu_dbus_sel[3] ),
    .CLK(net15),
    .Q(\u_arbiter.i_wb_cpu_rdt[3] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[60]  (.D(\u_scanchain_local.module_data_in[59] ),
    .SE(net554),
    .SI(\u_arbiter.o_wb_cpu_adr[22] ),
    .CLK(net22),
    .Q(\u_scanchain_local.module_data_in[60] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[61]  (.D(\u_scanchain_local.module_data_in[60] ),
    .SE(net555),
    .SI(\u_arbiter.o_wb_cpu_adr[23] ),
    .CLK(net23),
    .Q(\u_scanchain_local.module_data_in[61] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[62]  (.D(\u_scanchain_local.module_data_in[61] ),
    .SE(net555),
    .SI(\u_arbiter.o_wb_cpu_adr[24] ),
    .CLK(net22),
    .Q(\u_scanchain_local.module_data_in[62] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[63]  (.D(\u_scanchain_local.module_data_in[62] ),
    .SE(net556),
    .SI(\u_arbiter.o_wb_cpu_adr[25] ),
    .CLK(net24),
    .Q(\u_scanchain_local.module_data_in[63] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[64]  (.D(\u_scanchain_local.module_data_in[63] ),
    .SE(net554),
    .SI(\u_arbiter.o_wb_cpu_adr[26] ),
    .CLK(net23),
    .Q(\u_scanchain_local.module_data_in[64] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[65]  (.D(\u_scanchain_local.module_data_in[64] ),
    .SE(net554),
    .SI(\u_arbiter.o_wb_cpu_adr[27] ),
    .CLK(net22),
    .Q(\u_scanchain_local.module_data_in[65] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[66]  (.D(\u_scanchain_local.module_data_in[65] ),
    .SE(net554),
    .SI(\u_arbiter.o_wb_cpu_adr[28] ),
    .CLK(net22),
    .Q(\u_scanchain_local.module_data_in[66] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[67]  (.D(\u_scanchain_local.module_data_in[66] ),
    .SE(net554),
    .SI(\u_arbiter.o_wb_cpu_adr[29] ),
    .CLK(net22),
    .Q(\u_scanchain_local.module_data_in[67] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[68]  (.D(\u_scanchain_local.module_data_in[67] ),
    .SE(net559),
    .SI(\u_arbiter.o_wb_cpu_adr[30] ),
    .CLK(net27),
    .Q(\u_scanchain_local.module_data_in[68] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[69]  (.D(\u_scanchain_local.module_data_in[68] ),
    .SE(net559),
    .SI(\u_arbiter.o_wb_cpu_adr[31] ),
    .CLK(net27),
    .Q(\u_scanchain_local.module_data_in[69] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[6]  (.D(\u_arbiter.i_wb_cpu_rdt[3] ),
    .SE(net548),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[0] ),
    .CLK(net15),
    .Q(\u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[7]  (.D(\u_arbiter.i_wb_cpu_rdt[4] ),
    .SE(net548),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[1] ),
    .CLK(net15),
    .Q(\u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[8]  (.D(\u_arbiter.i_wb_cpu_rdt[5] ),
    .SE(net549),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[2] ),
    .CLK(net16),
    .Q(\u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[9]  (.D(\u_arbiter.i_wb_cpu_rdt[6] ),
    .SE(net544),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[3] ),
    .CLK(net12),
    .Q(\u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3892 ();
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input1 (.I(io_in[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input2 (.I(io_in[1]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input3 (.I(io_in[2]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input4 (.I(io_in[3]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input5 (.I(io_in[4]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output6 (.I(net6),
    .Z(io_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output7 (.I(net7),
    .Z(io_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout8 (.I(\u_arbiter.i_wb_cpu_ack ),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout9 (.I(net14),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout10 (.I(net11),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout11 (.I(net14),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout12 (.I(net14),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout13 (.I(net14),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout14 (.I(net19),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout15 (.I(net16),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout16 (.I(net18),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout17 (.I(net18),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout18 (.I(net19),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout19 (.I(net35),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout20 (.I(net25),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout21 (.I(net25),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout22 (.I(net24),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout23 (.I(net24),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout24 (.I(net25),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout25 (.I(net33),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout26 (.I(net28),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout27 (.I(net32),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout28 (.I(net32),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 fanout29 (.I(net31),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout30 (.I(net31),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout31 (.I(net32),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout32 (.I(net33),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout33 (.I(net34),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout34 (.I(net35),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout35 (.I(\u_scanchain_local.clk ),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout36 (.I(\u_arbiter.i_wb_cpu_dbus_dat[1] ),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout37 (.I(net43),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout38 (.I(net42),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout39 (.I(net42),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout40 (.I(net42),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout41 (.I(net42),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout42 (.I(net43),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout43 (.I(net50),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout44 (.I(net45),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout45 (.I(net49),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout46 (.I(net49),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout47 (.I(net48),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout48 (.I(net49),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout49 (.I(net50),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout50 (.I(net73),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout51 (.I(net55),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout52 (.I(net55),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout53 (.I(net55),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout54 (.I(net55),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout55 (.I(net62),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout56 (.I(net58),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout57 (.I(net58),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout58 (.I(net61),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout59 (.I(net61),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout60 (.I(net61),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout61 (.I(net62),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout62 (.I(net72),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout63 (.I(net65),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout64 (.I(net65),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout65 (.I(net71),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout66 (.I(net71),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout67 (.I(net70),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout68 (.I(net70),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout69 (.I(net70),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout70 (.I(net71),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout71 (.I(net72),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout72 (.I(net73),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout73 (.I(net109),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout74 (.I(net75),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout75 (.I(net78),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout76 (.I(net78),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout77 (.I(net78),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout78 (.I(net84),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 fanout79 (.I(net83),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout80 (.I(net83),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout81 (.I(net83),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout82 (.I(net83),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout83 (.I(net84),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout84 (.I(net92),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout85 (.I(net89),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout86 (.I(net89),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout87 (.I(net89),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout88 (.I(net89),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout89 (.I(net91),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout90 (.I(net91),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout91 (.I(net92),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout92 (.I(net108),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout93 (.I(net95),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout94 (.I(net95),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout95 (.I(net97),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout96 (.I(net97),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout97 (.I(net100),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout98 (.I(net99),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout99 (.I(net100),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout100 (.I(net107),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout101 (.I(net104),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout102 (.I(net104),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout103 (.I(net105),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout104 (.I(net105),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout105 (.I(net107),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout106 (.I(net107),
    .Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout107 (.I(net108),
    .Z(net107));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout108 (.I(net109),
    .Z(net108));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout109 (.I(net158),
    .Z(net109));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout110 (.I(net113),
    .Z(net110));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout111 (.I(net113),
    .Z(net111));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout112 (.I(net113),
    .Z(net112));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout113 (.I(net115),
    .Z(net113));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout114 (.I(net115),
    .Z(net114));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout115 (.I(net120),
    .Z(net115));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout116 (.I(net119),
    .Z(net116));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout117 (.I(net119),
    .Z(net117));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout118 (.I(net119),
    .Z(net118));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout119 (.I(net120),
    .Z(net119));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout120 (.I(net131),
    .Z(net120));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout121 (.I(net124),
    .Z(net121));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout122 (.I(net124),
    .Z(net122));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout123 (.I(net124),
    .Z(net123));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout124 (.I(net130),
    .Z(net124));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout125 (.I(net129),
    .Z(net125));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout126 (.I(net129),
    .Z(net126));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout127 (.I(net129),
    .Z(net127));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout128 (.I(net129),
    .Z(net128));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout129 (.I(net130),
    .Z(net129));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout130 (.I(net131),
    .Z(net130));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout131 (.I(net132),
    .Z(net131));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout132 (.I(net157),
    .Z(net132));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout133 (.I(net139),
    .Z(net133));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout134 (.I(net139),
    .Z(net134));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout135 (.I(net137),
    .Z(net135));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout136 (.I(net137),
    .Z(net136));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout137 (.I(net139),
    .Z(net137));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout138 (.I(net139),
    .Z(net138));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout139 (.I(net148),
    .Z(net139));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout140 (.I(net142),
    .Z(net140));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout141 (.I(net142),
    .Z(net141));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout142 (.I(net147),
    .Z(net142));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout143 (.I(net145),
    .Z(net143));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout144 (.I(net145),
    .Z(net144));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout145 (.I(net147),
    .Z(net145));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout146 (.I(net147),
    .Z(net146));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout147 (.I(net148),
    .Z(net147));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout148 (.I(net156),
    .Z(net148));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout149 (.I(net151),
    .Z(net149));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout150 (.I(net151),
    .Z(net150));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout151 (.I(net155),
    .Z(net151));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout152 (.I(net154),
    .Z(net152));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout153 (.I(net154),
    .Z(net153));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout154 (.I(net155),
    .Z(net154));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout155 (.I(net156),
    .Z(net155));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout156 (.I(net157),
    .Z(net156));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout157 (.I(net158),
    .Z(net157));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout158 (.I(net269),
    .Z(net158));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout159 (.I(net161),
    .Z(net159));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout160 (.I(net164),
    .Z(net160));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout161 (.I(net164),
    .Z(net161));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout162 (.I(net163),
    .Z(net162));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout163 (.I(net164),
    .Z(net163));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout164 (.I(net173),
    .Z(net164));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout165 (.I(net167),
    .Z(net165));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout166 (.I(net167),
    .Z(net166));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout167 (.I(net172),
    .Z(net167));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout168 (.I(net170),
    .Z(net168));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout169 (.I(net170),
    .Z(net169));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout170 (.I(net172),
    .Z(net170));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout171 (.I(net172),
    .Z(net171));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout172 (.I(net173),
    .Z(net172));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout173 (.I(net194),
    .Z(net173));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout174 (.I(net176),
    .Z(net174));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout175 (.I(net176),
    .Z(net175));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout176 (.I(net184),
    .Z(net176));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout177 (.I(net184),
    .Z(net177));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout178 (.I(net180),
    .Z(net178));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout179 (.I(net183),
    .Z(net179));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout180 (.I(net183),
    .Z(net180));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout181 (.I(net183),
    .Z(net181));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout182 (.I(net183),
    .Z(net182));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout183 (.I(net184),
    .Z(net183));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout184 (.I(net193),
    .Z(net184));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout185 (.I(net187),
    .Z(net185));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout186 (.I(net187),
    .Z(net186));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout187 (.I(net192),
    .Z(net187));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout188 (.I(net191),
    .Z(net188));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout189 (.I(net191),
    .Z(net189));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout190 (.I(net191),
    .Z(net190));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout191 (.I(net192),
    .Z(net191));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout192 (.I(net193),
    .Z(net192));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout193 (.I(net194),
    .Z(net193));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout194 (.I(net231),
    .Z(net194));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout195 (.I(net196),
    .Z(net195));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout196 (.I(net202),
    .Z(net196));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout197 (.I(net202),
    .Z(net197));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout198 (.I(net199),
    .Z(net198));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout199 (.I(net201),
    .Z(net199));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout200 (.I(net201),
    .Z(net200));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout201 (.I(net202),
    .Z(net201));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout202 (.I(net209),
    .Z(net202));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout203 (.I(net208),
    .Z(net203));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout204 (.I(net208),
    .Z(net204));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout205 (.I(net207),
    .Z(net205));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout206 (.I(net207),
    .Z(net206));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout207 (.I(net208),
    .Z(net207));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout208 (.I(net209),
    .Z(net208));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout209 (.I(net214),
    .Z(net209));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout210 (.I(net211),
    .Z(net210));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout211 (.I(net213),
    .Z(net211));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout212 (.I(net213),
    .Z(net212));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout213 (.I(net214),
    .Z(net213));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout214 (.I(net230),
    .Z(net214));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout215 (.I(net219),
    .Z(net215));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout216 (.I(net219),
    .Z(net216));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout217 (.I(net219),
    .Z(net217));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout218 (.I(net219),
    .Z(net218));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout219 (.I(net223),
    .Z(net219));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout220 (.I(net221),
    .Z(net220));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout221 (.I(net223),
    .Z(net221));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout222 (.I(net223),
    .Z(net222));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout223 (.I(net229),
    .Z(net223));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout224 (.I(net228),
    .Z(net224));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout225 (.I(net228),
    .Z(net225));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout226 (.I(net228),
    .Z(net226));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout227 (.I(net228),
    .Z(net227));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout228 (.I(net229),
    .Z(net228));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout229 (.I(net230),
    .Z(net229));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout230 (.I(net231),
    .Z(net230));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout231 (.I(net268),
    .Z(net231));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout232 (.I(net235),
    .Z(net232));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout233 (.I(net235),
    .Z(net233));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout234 (.I(net235),
    .Z(net234));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout235 (.I(net240),
    .Z(net235));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout236 (.I(net238),
    .Z(net236));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout237 (.I(net238),
    .Z(net237));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout238 (.I(net240),
    .Z(net238));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout239 (.I(net240),
    .Z(net239));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout240 (.I(net247),
    .Z(net240));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout241 (.I(net246),
    .Z(net241));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout242 (.I(net246),
    .Z(net242));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout243 (.I(net244),
    .Z(net243));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout244 (.I(net245),
    .Z(net244));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout245 (.I(net246),
    .Z(net245));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout246 (.I(net247),
    .Z(net246));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout247 (.I(net248),
    .Z(net247));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout248 (.I(net267),
    .Z(net248));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout249 (.I(net255),
    .Z(net249));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout250 (.I(net255),
    .Z(net250));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout251 (.I(net254),
    .Z(net251));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout252 (.I(net253),
    .Z(net252));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout253 (.I(net254),
    .Z(net253));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout254 (.I(net255),
    .Z(net254));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout255 (.I(net262),
    .Z(net255));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout256 (.I(net257),
    .Z(net256));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout257 (.I(net260),
    .Z(net257));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout258 (.I(net259),
    .Z(net258));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout259 (.I(net260),
    .Z(net259));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout260 (.I(net261),
    .Z(net260));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout261 (.I(net262),
    .Z(net261));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout262 (.I(net266),
    .Z(net262));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout263 (.I(net264),
    .Z(net263));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout264 (.I(net265),
    .Z(net264));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout265 (.I(net266),
    .Z(net265));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout266 (.I(net267),
    .Z(net266));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout267 (.I(net268),
    .Z(net267));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout268 (.I(net269),
    .Z(net268));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout269 (.I(net540),
    .Z(net269));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout270 (.I(net271),
    .Z(net270));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout271 (.I(net275),
    .Z(net271));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout272 (.I(net273),
    .Z(net272));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout273 (.I(net274),
    .Z(net273));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout274 (.I(net275),
    .Z(net274));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout275 (.I(net281),
    .Z(net275));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout276 (.I(net280),
    .Z(net276));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout277 (.I(net280),
    .Z(net277));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout278 (.I(net279),
    .Z(net278));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout279 (.I(net280),
    .Z(net279));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout280 (.I(net281),
    .Z(net280));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout281 (.I(net290),
    .Z(net281));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout282 (.I(net283),
    .Z(net282));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout283 (.I(net284),
    .Z(net283));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout284 (.I(net285),
    .Z(net284));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout285 (.I(net289),
    .Z(net285));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout286 (.I(net288),
    .Z(net286));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout287 (.I(net288),
    .Z(net287));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout288 (.I(net289),
    .Z(net288));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout289 (.I(net290),
    .Z(net289));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout290 (.I(net306),
    .Z(net290));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout291 (.I(net294),
    .Z(net291));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout292 (.I(net294),
    .Z(net292));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout293 (.I(net294),
    .Z(net293));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout294 (.I(net298),
    .Z(net294));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout295 (.I(net298),
    .Z(net295));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout296 (.I(net297),
    .Z(net296));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout297 (.I(net298),
    .Z(net297));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout298 (.I(net305),
    .Z(net298));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 fanout299 (.I(net304),
    .Z(net299));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout300 (.I(net304),
    .Z(net300));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout301 (.I(net303),
    .Z(net301));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout302 (.I(net303),
    .Z(net302));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout303 (.I(net304),
    .Z(net303));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout304 (.I(net305),
    .Z(net304));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout305 (.I(net306),
    .Z(net305));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout306 (.I(net338),
    .Z(net306));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout307 (.I(net311),
    .Z(net307));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout308 (.I(net311),
    .Z(net308));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout309 (.I(net310),
    .Z(net309));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout310 (.I(net311),
    .Z(net310));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout311 (.I(net315),
    .Z(net311));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout312 (.I(net315),
    .Z(net312));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout313 (.I(net314),
    .Z(net313));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout314 (.I(net315),
    .Z(net314));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout315 (.I(net323),
    .Z(net315));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout316 (.I(net317),
    .Z(net316));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout317 (.I(net322),
    .Z(net317));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout318 (.I(net322),
    .Z(net318));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout319 (.I(net320),
    .Z(net319));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout320 (.I(net322),
    .Z(net320));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout321 (.I(net322),
    .Z(net321));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout322 (.I(net323),
    .Z(net322));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout323 (.I(net337),
    .Z(net323));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout324 (.I(net325),
    .Z(net324));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout325 (.I(net328),
    .Z(net325));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 fanout326 (.I(net328),
    .Z(net326));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout327 (.I(net328),
    .Z(net327));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout328 (.I(net336),
    .Z(net328));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout329 (.I(net332),
    .Z(net329));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout330 (.I(net332),
    .Z(net330));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout331 (.I(net332),
    .Z(net331));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout332 (.I(net335),
    .Z(net332));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout333 (.I(net334),
    .Z(net333));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout334 (.I(net335),
    .Z(net334));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout335 (.I(net336),
    .Z(net335));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout336 (.I(net337),
    .Z(net336));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout337 (.I(net338),
    .Z(net337));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout338 (.I(net395),
    .Z(net338));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout339 (.I(net340),
    .Z(net339));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout340 (.I(net345),
    .Z(net340));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout341 (.I(net344),
    .Z(net341));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout342 (.I(net344),
    .Z(net342));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout343 (.I(net344),
    .Z(net343));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout344 (.I(net345),
    .Z(net344));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout345 (.I(net356),
    .Z(net345));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout346 (.I(net349),
    .Z(net346));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 fanout347 (.I(net349),
    .Z(net347));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout348 (.I(net349),
    .Z(net348));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout349 (.I(net355),
    .Z(net349));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout350 (.I(net354),
    .Z(net350));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout351 (.I(net354),
    .Z(net351));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout352 (.I(net354),
    .Z(net352));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout353 (.I(net354),
    .Z(net353));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout354 (.I(net355),
    .Z(net354));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout355 (.I(net356),
    .Z(net355));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout356 (.I(net367),
    .Z(net356));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout357 (.I(net366),
    .Z(net357));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout358 (.I(net359),
    .Z(net358));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout359 (.I(net366),
    .Z(net359));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout360 (.I(net362),
    .Z(net360));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout361 (.I(net362),
    .Z(net361));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout362 (.I(net365),
    .Z(net362));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout363 (.I(net365),
    .Z(net363));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout364 (.I(net365),
    .Z(net364));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout365 (.I(net366),
    .Z(net365));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout366 (.I(net367),
    .Z(net366));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout367 (.I(net394),
    .Z(net367));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout368 (.I(net372),
    .Z(net368));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout369 (.I(net372),
    .Z(net369));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout370 (.I(net372),
    .Z(net370));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout371 (.I(net372),
    .Z(net371));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout372 (.I(net375),
    .Z(net372));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout373 (.I(net374),
    .Z(net373));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout374 (.I(net375),
    .Z(net374));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout375 (.I(net382),
    .Z(net375));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout376 (.I(net381),
    .Z(net376));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout377 (.I(net381),
    .Z(net377));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout378 (.I(net380),
    .Z(net378));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout379 (.I(net380),
    .Z(net379));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout380 (.I(net381),
    .Z(net380));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout381 (.I(net382),
    .Z(net381));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout382 (.I(net393),
    .Z(net382));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout383 (.I(net384),
    .Z(net383));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout384 (.I(net385),
    .Z(net384));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout385 (.I(net388),
    .Z(net385));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout386 (.I(net387),
    .Z(net386));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 fanout387 (.I(net388),
    .Z(net387));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout388 (.I(net392),
    .Z(net388));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout389 (.I(net391),
    .Z(net389));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout390 (.I(net391),
    .Z(net390));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout391 (.I(net392),
    .Z(net391));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout392 (.I(net393),
    .Z(net392));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout393 (.I(net394),
    .Z(net393));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout394 (.I(net395),
    .Z(net394));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout395 (.I(net539),
    .Z(net395));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout396 (.I(net397),
    .Z(net396));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout397 (.I(net399),
    .Z(net397));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout398 (.I(net399),
    .Z(net398));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout399 (.I(net402),
    .Z(net399));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout400 (.I(net402),
    .Z(net400));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout401 (.I(net402),
    .Z(net401));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout402 (.I(net414),
    .Z(net402));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout403 (.I(net407),
    .Z(net403));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout404 (.I(net407),
    .Z(net404));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout405 (.I(net406),
    .Z(net405));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout406 (.I(net407),
    .Z(net406));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout407 (.I(net413),
    .Z(net407));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout408 (.I(net412),
    .Z(net408));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout409 (.I(net412),
    .Z(net409));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout410 (.I(net412),
    .Z(net410));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout411 (.I(net412),
    .Z(net411));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout412 (.I(net413),
    .Z(net412));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout413 (.I(net414),
    .Z(net413));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout414 (.I(net435),
    .Z(net414));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout415 (.I(net417),
    .Z(net415));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout416 (.I(net417),
    .Z(net416));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout417 (.I(net424),
    .Z(net417));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout418 (.I(net424),
    .Z(net418));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout419 (.I(net423),
    .Z(net419));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout420 (.I(net423),
    .Z(net420));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout421 (.I(net423),
    .Z(net421));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout422 (.I(net423),
    .Z(net422));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout423 (.I(net424),
    .Z(net423));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout424 (.I(net434),
    .Z(net424));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout425 (.I(net429),
    .Z(net425));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout426 (.I(net429),
    .Z(net426));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout427 (.I(net428),
    .Z(net427));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout428 (.I(net429),
    .Z(net428));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout429 (.I(net433),
    .Z(net429));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout430 (.I(net431),
    .Z(net430));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout431 (.I(net433),
    .Z(net431));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout432 (.I(net433),
    .Z(net432));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout433 (.I(net434),
    .Z(net433));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout434 (.I(net435),
    .Z(net434));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout435 (.I(net476),
    .Z(net435));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout436 (.I(net442),
    .Z(net436));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout437 (.I(net442),
    .Z(net437));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout438 (.I(net440),
    .Z(net438));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout439 (.I(net440),
    .Z(net439));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout440 (.I(net442),
    .Z(net440));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout441 (.I(net442),
    .Z(net441));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout442 (.I(net449),
    .Z(net442));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout443 (.I(net444),
    .Z(net443));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout444 (.I(net447),
    .Z(net444));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout445 (.I(net446),
    .Z(net445));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout446 (.I(net447),
    .Z(net446));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout447 (.I(net448),
    .Z(net447));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout448 (.I(net449),
    .Z(net448));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout449 (.I(net475),
    .Z(net449));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout450 (.I(net452),
    .Z(net450));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout451 (.I(net452),
    .Z(net451));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout452 (.I(net455),
    .Z(net452));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout453 (.I(net455),
    .Z(net453));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout454 (.I(net455),
    .Z(net454));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout455 (.I(net460),
    .Z(net455));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout456 (.I(net457),
    .Z(net456));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout457 (.I(net459),
    .Z(net457));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout458 (.I(net459),
    .Z(net458));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout459 (.I(net460),
    .Z(net459));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout460 (.I(net474),
    .Z(net460));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout461 (.I(net467),
    .Z(net461));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout462 (.I(net467),
    .Z(net462));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout463 (.I(net466),
    .Z(net463));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout464 (.I(net466),
    .Z(net464));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout465 (.I(net467),
    .Z(net465));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout466 (.I(net467),
    .Z(net466));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout467 (.I(net473),
    .Z(net467));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout468 (.I(net469),
    .Z(net468));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout469 (.I(net472),
    .Z(net469));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout470 (.I(net471),
    .Z(net470));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout471 (.I(net472),
    .Z(net471));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout472 (.I(net473),
    .Z(net472));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout473 (.I(net474),
    .Z(net473));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout474 (.I(net475),
    .Z(net474));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout475 (.I(net476),
    .Z(net475));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout476 (.I(net538),
    .Z(net476));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout477 (.I(net484),
    .Z(net477));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout478 (.I(net484),
    .Z(net478));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout479 (.I(net483),
    .Z(net479));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout480 (.I(net483),
    .Z(net480));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout481 (.I(net483),
    .Z(net481));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout482 (.I(net483),
    .Z(net482));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout483 (.I(net484),
    .Z(net483));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout484 (.I(net494),
    .Z(net484));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout485 (.I(net487),
    .Z(net485));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout486 (.I(net487),
    .Z(net486));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout487 (.I(net489),
    .Z(net487));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout488 (.I(net489),
    .Z(net488));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout489 (.I(net493),
    .Z(net489));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout490 (.I(net492),
    .Z(net490));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout491 (.I(net492),
    .Z(net491));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout492 (.I(net493),
    .Z(net492));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout493 (.I(net494),
    .Z(net493));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout494 (.I(net507),
    .Z(net494));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout495 (.I(net499),
    .Z(net495));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout496 (.I(net499),
    .Z(net496));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 fanout497 (.I(net499),
    .Z(net497));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout498 (.I(net499),
    .Z(net498));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout499 (.I(net506),
    .Z(net499));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout500 (.I(net502),
    .Z(net500));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout501 (.I(net502),
    .Z(net501));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout502 (.I(net505),
    .Z(net502));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout503 (.I(net505),
    .Z(net503));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout504 (.I(net505),
    .Z(net504));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout505 (.I(net506),
    .Z(net505));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout506 (.I(net507),
    .Z(net506));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout507 (.I(net537),
    .Z(net507));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout508 (.I(net509),
    .Z(net508));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout509 (.I(net510),
    .Z(net509));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout510 (.I(net511),
    .Z(net510));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout511 (.I(net515),
    .Z(net511));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout512 (.I(net514),
    .Z(net512));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout513 (.I(net514),
    .Z(net513));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout514 (.I(net515),
    .Z(net514));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout515 (.I(net522),
    .Z(net515));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout516 (.I(net520),
    .Z(net516));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout517 (.I(net520),
    .Z(net517));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout518 (.I(net519),
    .Z(net518));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout519 (.I(net520),
    .Z(net519));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout520 (.I(net521),
    .Z(net520));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout521 (.I(net522),
    .Z(net521));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout522 (.I(net536),
    .Z(net522));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout523 (.I(net527),
    .Z(net523));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout524 (.I(net527),
    .Z(net524));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout525 (.I(net527),
    .Z(net525));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout526 (.I(net527),
    .Z(net526));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout527 (.I(net535),
    .Z(net527));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout528 (.I(net530),
    .Z(net528));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout529 (.I(net530),
    .Z(net529));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout530 (.I(net534),
    .Z(net530));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout531 (.I(net534),
    .Z(net531));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout532 (.I(net534),
    .Z(net532));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout533 (.I(net534),
    .Z(net533));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout534 (.I(net535),
    .Z(net534));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout535 (.I(net536),
    .Z(net535));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout536 (.I(net537),
    .Z(net536));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout537 (.I(net538),
    .Z(net537));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout538 (.I(net539),
    .Z(net538));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout539 (.I(net540),
    .Z(net539));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout540 (.I(net5),
    .Z(net540));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout541 (.I(net543),
    .Z(net541));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout542 (.I(net546),
    .Z(net542));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout543 (.I(net546),
    .Z(net543));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout544 (.I(net546),
    .Z(net544));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout545 (.I(net546),
    .Z(net545));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout546 (.I(net551),
    .Z(net546));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout547 (.I(net550),
    .Z(net547));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout548 (.I(net549),
    .Z(net548));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout549 (.I(net550),
    .Z(net549));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout550 (.I(net551),
    .Z(net550));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout551 (.I(net565),
    .Z(net551));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout552 (.I(net557),
    .Z(net552));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout553 (.I(net557),
    .Z(net553));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout554 (.I(net556),
    .Z(net554));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout555 (.I(net556),
    .Z(net555));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout556 (.I(net557),
    .Z(net556));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout557 (.I(net564),
    .Z(net557));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout558 (.I(net560),
    .Z(net558));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout559 (.I(net563),
    .Z(net559));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout560 (.I(net563),
    .Z(net560));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout561 (.I(net562),
    .Z(net561));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout562 (.I(net563),
    .Z(net562));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout563 (.I(net564),
    .Z(net563));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout564 (.I(net565),
    .Z(net564));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout565 (.I(net4),
    .Z(net565));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06410__A1 (.I(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06298__A1 (.I(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06142__A1 (.I(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05778__A3 (.I(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06525__I (.I(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06309__I (.I(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06140__I (.I(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06064__I (.I(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05776__I (.I(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06856__C (.I(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06768__C (.I(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06680__C (.I(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06167__I (.I(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05777__I (.I(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06475__C (.I(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06361__C (.I(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06245__C (.I(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06029__C (.I(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05778__A4 (.I(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07072__A1 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07070__A1 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07067__A1 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07065__A1 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05781__I (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10286__A1 (.I(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07109__A1 (.I(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07103__A1 (.I(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06972__A1 (.I(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05786__A1 (.I(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09145__A1 (.I(_01432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09129__I (.I(_01432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05803__A1 (.I(_01432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05784__A1 (.I(_01432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09740__A2 (.I(_01433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07694__A2 (.I(_01433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05788__A2 (.I(_01433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05785__I (.I(_01433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07089__A2 (.I(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05945__S (.I(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05826__A1 (.I(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05802__A1 (.I(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05786__A2 (.I(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09688__I (.I(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09676__S (.I(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09674__S (.I(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07691__I (.I(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05791__I (.I(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09724__A1 (.I(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09715__A1 (.I(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09677__S (.I(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09675__S (.I(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05792__I (.I(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10026__A1 (.I(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09994__A1 (.I(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09895__S (.I(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09685__A1 (.I(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05794__I (.I(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10087__S (.I(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09936__S (.I(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09893__S (.I(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05799__I (.I(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05795__I (.I(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10574__A1 (.I(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10001__A1 (.I(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09989__A1 (.I(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09969__A1 (.I(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05798__A1 (.I(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10072__S (.I(_01446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09984__S (.I(_01446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09952__S (.I(_01446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09859__S (.I(_01446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05800__I (.I(_01446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10118__S (.I(_01447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10011__S (.I(_01447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09843__S (.I(_01447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05814__A1 (.I(_01447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05801__A1 (.I(_01447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09527__A2 (.I(_01450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07711__A2 (.I(_01450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05804__I (.I(_01450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05914__I (.I(_01451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05879__I (.I(_01451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05855__I (.I(_01451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05809__I (.I(_01451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05805__I (.I(_01451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05871__I (.I(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05851__I (.I(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05841__I (.I(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05816__I (.I(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05806__I (.I(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05911__A1 (.I(_01453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05866__A2 (.I(_01453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05844__A2 (.I(_01453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05812__A2 (.I(_01453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05807__A2 (.I(_01453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05896__I (.I(_01455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05868__B (.I(_01455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05848__B (.I(_01455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05832__I (.I(_01455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05810__I (.I(_01455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07087__B (.I(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05831__A1 (.I(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05823__A1 (.I(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05818__A1 (.I(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05813__A1 (.I(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05838__A2 (.I(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05830__A2 (.I(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05827__A2 (.I(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05822__A2 (.I(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05817__A2 (.I(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10298__A1 (.I(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10295__B2 (.I(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05825__A2 (.I(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05824__A1 (.I(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05821__A1 (.I(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05834__A4 (.I(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05825__A3 (.I(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05824__A2 (.I(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05821__A2 (.I(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05895__A1 (.I(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05884__A1 (.I(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05861__A1 (.I(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05843__A1 (.I(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05839__A1 (.I(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05899__A2 (.I(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05894__A2 (.I(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05883__A2 (.I(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05860__A2 (.I(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05842__A2 (.I(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05941__A1 (.I(_01489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05937__A1 (.I(_01489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05933__A1 (.I(_01489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05865__A1 (.I(_01489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05857__A1 (.I(_01489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05940__A2 (.I(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05936__A2 (.I(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05875__A2 (.I(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05864__A2 (.I(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05856__A2 (.I(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05906__A1 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05892__A1 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05888__A1 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05881__A1 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05876__A1 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05910__A2 (.I(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05905__A2 (.I(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05891__A2 (.I(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05887__A2 (.I(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05880__A2 (.I(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05902__A4 (.I(_01516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05890__A2 (.I(_01516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05889__A2 (.I(_01516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05888__A2 (.I(_01516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05929__A1 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05924__A1 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05920__A1 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05916__A1 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05900__A1 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05926__A4 (.I(_01535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05921__A3 (.I(_01535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05917__A2 (.I(_01535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05913__A2 (.I(_01535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05911__A3 (.I(_01535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10343__A1 (.I(_01537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10340__B2 (.I(_01537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05921__A2 (.I(_01537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05917__A1 (.I(_01537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05913__A1 (.I(_01537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05932__A2 (.I(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05928__A2 (.I(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05923__A2 (.I(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05919__A2 (.I(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05915__A2 (.I(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05943__A2 (.I(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05939__A2 (.I(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06905__A1 (.I(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06411__I (.I(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06143__I (.I(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05949__I (.I(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06085__I (.I(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06054__I (.I(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05978__I (.I(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05951__I (.I(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06445__I (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06213__I (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06202__I (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06066__I (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05952__I (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06914__A1 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06453__A1 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06340__A1 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06224__A1 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05962__A1 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06087__I (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06056__I (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06021__I (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06003__I (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05955__I (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06432__I (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06306__I (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06175__I (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06162__I (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05956__I (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06470__I (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06233__I (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06014__I (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05974__I (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05957__I (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06566__S0 (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06452__S0 (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06339__S0 (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06223__S0 (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05961__S0 (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06171__I (.I(_01575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06024__I (.I(_01575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05998__I (.I(_01575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05967__I (.I(_01575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05959__I (.I(_01575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06872__S1 (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06784__S1 (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06222__I (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05975__I (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05960__I (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06843__S1 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06755__S1 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06667__S1 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06579__S1 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05961__S1 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05962__A2 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06835__A1 (.I(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06456__A1 (.I(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06342__A1 (.I(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06227__A1 (.I(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05972__A1 (.I(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06195__I (.I(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06068__I (.I(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06033__I (.I(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05995__I (.I(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05965__I (.I(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06460__I (.I(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06321__S0 (.I(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06187__S0 (.I(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05981__I (.I(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05966__I (.I(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06568__S0 (.I(_01583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06454__S0 (.I(_01583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06341__S0 (.I(_01583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06226__S0 (.I(_01583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05969__S0 (.I(_01583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06425__I (.I(_01584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06225__I (.I(_01584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06182__I (.I(_01584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05982__I (.I(_01584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05968__I (.I(_01584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06836__S1 (.I(_01585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06748__S1 (.I(_01585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06660__S1 (.I(_01585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06572__S1 (.I(_01585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05969__S1 (.I(_01585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05972__A2 (.I(_01586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06871__B (.I(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06783__B (.I(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06695__B (.I(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06243__I (.I(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05971__I (.I(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06846__B (.I(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06758__B (.I(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06342__B (.I(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06227__B (.I(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05972__B (.I(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06844__A1 (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06756__A1 (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06668__A1 (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06229__A1 (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05977__A1 (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06830__S0 (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06742__S0 (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06654__S0 (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06228__S0 (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05976__S0 (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06830__S1 (.I(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06742__S1 (.I(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06345__S1 (.I(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06228__S1 (.I(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05976__S1 (.I(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05977__A2 (.I(_01593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06389__I (.I(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06111__I (.I(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06103__I (.I(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06039__I (.I(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05979__I (.I(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06467__I (.I(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06241__I (.I(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06020__I (.I(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06002__I (.I(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05980__I (.I(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06573__A1 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06462__A1 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06348__A1 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06231__A1 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05987__A1 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06841__S0 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06753__S0 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06347__S0 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06230__S0 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05983__S0 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06841__S1 (.I(_01599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06461__S1 (.I(_01599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06347__S1 (.I(_01599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06230__S1 (.I(_01599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05983__S1 (.I(_01599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05987__A2 (.I(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06251__I (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06045__I (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06010__I (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05985__I (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06851__B (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06763__B (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06355__I (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06206__I (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05986__I (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06842__B (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06462__B (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06348__B (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06231__B (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05987__B (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06284__I (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06116__I (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06094__I (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05989__I (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06876__C (.I(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06788__C (.I(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06435__I (.I(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06190__I (.I(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05990__I (.I(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06574__C (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06463__C (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06349__C (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06232__C (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05991__C (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06097__A2 (.I(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06536__I (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06373__I (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06134__I (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06074__I (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05993__I (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06860__A1 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06464__I (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06331__I (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06208__I (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05994__I (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06912__A1 (.I(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06824__A1 (.I(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06352__A1 (.I(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06235__A1 (.I(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06001__A1 (.I(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06318__I (.I(_01612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06181__I (.I(_01612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06170__I (.I(_01612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06145__I (.I(_01612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05996__I (.I(_01612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06446__I (.I(_01613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06214__I (.I(_01613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06209__I (.I(_01613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06203__I (.I(_01613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05997__I (.I(_01613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06911__S0 (.I(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06823__S0 (.I(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06735__S0 (.I(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06647__S0 (.I(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06000__S0 (.I(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06868__S1 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06780__S1 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06692__S1 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06350__I (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05999__I (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06911__S1 (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06823__S1 (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06735__S1 (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06234__S1 (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06000__S1 (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06846__A1 (.I(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06758__A1 (.I(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06356__A1 (.I(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06238__A1 (.I(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06012__A1 (.I(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06390__I (.I(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06104__I (.I(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06075__I (.I(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06040__I (.I(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06004__I (.I(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06394__S0 (.I(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06280__S0 (.I(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06236__I (.I(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06109__S0 (.I(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06005__I (.I(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06845__S0 (.I(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06757__S0 (.I(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06669__S0 (.I(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06581__S0 (.I(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06009__S0 (.I(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06859__S1 (.I(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06771__S1 (.I(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06353__I (.I(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06105__S1 (.I(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06008__I (.I(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06845__S1 (.I(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06757__S1 (.I(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06669__S1 (.I(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06237__S1 (.I(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06009__S1 (.I(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06012__A2 (.I(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06539__I (.I(_01627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06316__I (.I(_01627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06178__I (.I(_01627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06165__I (.I(_01627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06011__I (.I(_01627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06910__B (.I(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06822__B (.I(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06734__B (.I(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06238__B (.I(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06012__B (.I(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06580__A1 (.I(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06472__A1 (.I(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06358__A1 (.I(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06240__A1 (.I(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06019__A1 (.I(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06839__S0 (.I(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06751__S0 (.I(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06357__S0 (.I(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06239__S0 (.I(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06018__S0 (.I(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06537__I (.I(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06314__I (.I(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06176__I (.I(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06163__I (.I(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06016__I (.I(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06852__S1 (.I(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06764__S1 (.I(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06676__S1 (.I(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06109__S1 (.I(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06017__I (.I(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06839__S1 (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06471__S1 (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06357__S1 (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06239__S1 (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06018__S1 (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06019__A2 (.I(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06831__A1 (.I(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06743__A1 (.I(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06655__A1 (.I(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06567__A1 (.I(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06028__A1 (.I(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06508__I (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06481__I (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06386__I (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06099__I (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06022__I (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06868__S0 (.I(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06366__S0 (.I(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06253__S0 (.I(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06052__S0 (.I(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06023__I (.I(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06834__S0 (.I(_01640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06473__S0 (.I(_01640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06359__S0 (.I(_01640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06242__S0 (.I(_01640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06026__S0 (.I(_01640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06512__S1 (.I(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06396__S1 (.I(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06282__S1 (.I(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06113__S1 (.I(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06025__I (.I(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06581__S1 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06473__S1 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06359__S1 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06242__S1 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06026__S1 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06028__A2 (.I(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06914__B (.I(_01644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06826__B (.I(_01644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06738__B (.I(_01644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06650__B (.I(_01644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06028__B (.I(_01644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06097__A3 (.I(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06886__A1 (.I(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06798__A1 (.I(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06710__A1 (.I(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06622__A1 (.I(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06096__A1 (.I(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06399__I (.I(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06144__I (.I(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06118__I (.I(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06080__I (.I(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06032__I (.I(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06878__A1 (.I(_01649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06477__A1 (.I(_01649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06363__A1 (.I(_01649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06249__A1 (.I(_01649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06038__A1 (.I(_01649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06519__I (.I(_01650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06247__I (.I(_01650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06130__I (.I(_01650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06081__I (.I(_01650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06034__I (.I(_01650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06891__S0 (.I(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06803__S0 (.I(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06715__S0 (.I(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06627__S0 (.I(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06037__S0 (.I(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06418__I (.I(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06292__I (.I(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06157__I (.I(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06131__I (.I(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06036__I (.I(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06891__S1 (.I(_01653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06476__S1 (.I(_01653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06362__S1 (.I(_01653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06248__S1 (.I(_01653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06037__S1 (.I(_01653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06065__A1 (.I(_01655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06871__A1 (.I(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06480__A1 (.I(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06365__A1 (.I(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06252__A1 (.I(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06047__A1 (.I(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06870__S0 (.I(_01657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06479__S0 (.I(_01657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06364__S0 (.I(_01657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06250__S0 (.I(_01657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06044__S0 (.I(_01657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07279__A1 (.I(_01658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07139__A1 (.I(_01658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06089__I (.I(_01658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06058__I (.I(_01658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06042__I (.I(_01658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06478__I (.I(_01659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06276__I (.I(_01659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06263__I (.I(_01659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06076__I (.I(_01659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06043__I (.I(_01659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06870__S1 (.I(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06782__S1 (.I(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06364__S1 (.I(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06250__S1 (.I(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06044__S1 (.I(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06047__A2 (.I(_01661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06381__I (.I(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06138__I (.I(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06114__I (.I(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06092__I (.I(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06046__I (.I(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06875__B (.I(_01663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06787__B (.I(_01663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06699__B (.I(_01663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06611__B (.I(_01663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06047__B (.I(_01663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06503__I (.I(_01665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06266__I (.I(_01665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06108__I (.I(_01665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06098__I (.I(_01665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06049__I (.I(_01665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06495__I (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06279__I (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06100__I (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06082__I (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06051__I (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06065__B1 (.I(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06484__I (.I(_01671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06288__I (.I(_01671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06149__I (.I(_01671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06123__I (.I(_01671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06055__I (.I(_01671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06880__A1 (.I(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06792__A1 (.I(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06369__A1 (.I(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06258__A1 (.I(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06063__A1 (.I(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06511__I (.I(_01673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06255__I (.I(_01673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06124__I (.I(_01673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06112__I (.I(_01673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06057__I (.I(_01673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06879__S0 (.I(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06791__S0 (.I(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06703__S0 (.I(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06615__S0 (.I(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06060__S0 (.I(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06485__I (.I(_01675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06289__I (.I(_01675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06151__I (.I(_01675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06125__I (.I(_01675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06059__I (.I(_01675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06879__S1 (.I(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06791__S1 (.I(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06368__S1 (.I(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06256__S1 (.I(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06060__S1 (.I(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06416__I (.I(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06257__I (.I(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06127__I (.I(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06078__I (.I(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06062__I (.I(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06880__B (.I(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06792__B (.I(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06704__B (.I(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06616__B (.I(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06063__B (.I(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06065__B2 (.I(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06096__A2 (.I(_01682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06424__I (.I(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06260__I (.I(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06180__I (.I(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06169__I (.I(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06067__I (.I(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06901__A1 (.I(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06813__A1 (.I(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06725__A1 (.I(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06637__A1 (.I(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06073__A1 (.I(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06528__I (.I(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06400__I (.I(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06156__I (.I(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06119__I (.I(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06069__I (.I(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06593__S0 (.I(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06490__S0 (.I(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06371__S0 (.I(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06261__S0 (.I(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06072__S0 (.I(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06489__I (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06299__I (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06146__I (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06120__I (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06071__I (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06887__S1 (.I(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06799__S1 (.I(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06371__S1 (.I(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06261__S1 (.I(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06072__S1 (.I(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06095__A1 (.I(_01690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06884__A1 (.I(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06796__A1 (.I(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06708__A1 (.I(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06265__A1 (.I(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06079__A1 (.I(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06595__S0 (.I(_01692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06492__S0 (.I(_01692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06374__S0 (.I(_01692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06264__S0 (.I(_01692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06077__S0 (.I(_01692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06874__S1 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06786__S1 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06698__S1 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06610__S1 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06077__S1 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06079__A2 (.I(_01694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06855__B (.I(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06767__B (.I(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06375__B (.I(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06265__B (.I(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06079__B (.I(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06881__S1 (.I(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06793__S1 (.I(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06376__S1 (.I(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06267__S1 (.I(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06083__S1 (.I(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06084__A2 (.I(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06095__B1 (.I(_01701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06533__I (.I(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06378__I (.I(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06155__I (.I(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06129__I (.I(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06086__I (.I(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06882__A1 (.I(_01703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06794__A1 (.I(_01703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06706__A1 (.I(_01703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06270__A1 (.I(_01703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06093__A1 (.I(_01703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06522__I (.I(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06414__I (.I(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06150__I (.I(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06135__I (.I(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06088__I (.I(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06599__S0 (.I(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06498__S0 (.I(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06380__S0 (.I(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06269__S0 (.I(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06091__S0 (.I(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06379__I (.I(_01706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06198__I (.I(_01706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06186__I (.I(_01706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06136__I (.I(_01706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06090__I (.I(_01706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06883__S1 (.I(_01707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06795__S1 (.I(_01707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06707__S1 (.I(_01707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06269__S1 (.I(_01707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06091__S1 (.I(_01707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06093__A2 (.I(_01708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06884__B (.I(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06796__B (.I(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06708__B (.I(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06270__B (.I(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06093__B (.I(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06095__B2 (.I(_01710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06904__C (.I(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06500__C (.I(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06383__C (.I(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06271__C (.I(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06095__C (.I(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06097__B (.I(_01713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06862__A1 (.I(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06774__A1 (.I(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06388__A1 (.I(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06275__A1 (.I(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06102__A1 (.I(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06861__S0 (.I(_01716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06773__S0 (.I(_01716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06685__S0 (.I(_01716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06274__S0 (.I(_01716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06101__S0 (.I(_01716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06604__S1 (.I(_01717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06504__S1 (.I(_01717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06387__S1 (.I(_01717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06274__S1 (.I(_01717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06101__S1 (.I(_01717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06117__A1 (.I(_01719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06859__S0 (.I(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06771__S0 (.I(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06683__S0 (.I(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06277__S0 (.I(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06105__S0 (.I(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06107__A2 (.I(_01722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06117__A2 (.I(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06853__A1 (.I(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06765__A1 (.I(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06677__A1 (.I(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06281__A1 (.I(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06110__A1 (.I(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06854__S0 (.I(_01729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06766__S0 (.I(_01729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06396__S0 (.I(_01729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06282__S0 (.I(_01729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06113__S0 (.I(_01729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06115__A2 (.I(_01730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06864__B (.I(_01731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06513__B (.I(_01731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06397__B (.I(_01731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06283__B (.I(_01731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06115__B (.I(_01731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06865__C (.I(_01733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06777__C (.I(_01733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06689__C (.I(_01733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06601__C (.I(_01733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06117__C (.I(_01733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06142__A2 (.I(_01734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06888__A1 (.I(_01735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06800__A1 (.I(_01735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06712__A1 (.I(_01735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06287__A1 (.I(_01735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06122__A1 (.I(_01735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06857__S0 (.I(_01736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06769__S0 (.I(_01736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06681__S0 (.I(_01736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06286__S0 (.I(_01736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06121__S0 (.I(_01736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06613__S1 (.I(_01737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06515__S1 (.I(_01737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06401__S1 (.I(_01737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06286__S1 (.I(_01737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06121__S1 (.I(_01737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06122__A2 (.I(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06890__A1 (.I(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06802__A1 (.I(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06714__A1 (.I(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06626__A1 (.I(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06128__A1 (.I(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06889__S0 (.I(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06517__S0 (.I(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06403__S0 (.I(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06290__S0 (.I(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06126__S0 (.I(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06889__S1 (.I(_01742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06801__S1 (.I(_01742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06713__S1 (.I(_01742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06625__S1 (.I(_01742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06126__S1 (.I(_01742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06128__A2 (.I(_01743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06890__B (.I(_01744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06518__B (.I(_01744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06404__B (.I(_01744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06291__B (.I(_01744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06128__B (.I(_01744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06618__A1 (.I(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06521__A1 (.I(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06406__A1 (.I(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06294__A1 (.I(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06133__A1 (.I(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06848__S0 (.I(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06760__S0 (.I(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06405__S0 (.I(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06293__S0 (.I(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06132__S0 (.I(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06848__S1 (.I(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06760__S1 (.I(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06672__S1 (.I(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06584__S1 (.I(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06132__S1 (.I(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06133__A2 (.I(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06893__S0 (.I(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06805__S0 (.I(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06407__S0 (.I(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06295__S0 (.I(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06137__S0 (.I(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06141__B2 (.I(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06895__C (.I(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06807__C (.I(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06409__C (.I(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06297__C (.I(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06141__C (.I(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06142__A3 (.I(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06194__A1 (.I(_01759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06624__A1 (.I(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06530__A1 (.I(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06413__A1 (.I(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06301__A1 (.I(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06148__A1 (.I(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06900__S0 (.I(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06812__S0 (.I(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06412__S0 (.I(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06300__S0 (.I(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06147__S0 (.I(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06900__S1 (.I(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06812__S1 (.I(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06724__S1 (.I(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06636__S1 (.I(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06147__S1 (.I(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06168__A1 (.I(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06864__A1 (.I(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06532__A1 (.I(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06417__A1 (.I(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06303__A1 (.I(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06154__A1 (.I(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06863__S0 (.I(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06775__S0 (.I(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06687__S0 (.I(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06302__S0 (.I(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06152__S0 (.I(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06863__S1 (.I(_01768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06531__S1 (.I(_01768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06415__S1 (.I(_01768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06302__S1 (.I(_01768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06152__S1 (.I(_01768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06903__B (.I(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06815__B (.I(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06727__B (.I(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06303__B (.I(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06154__B (.I(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06168__A2 (.I(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06858__A1 (.I(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06770__A1 (.I(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06420__A1 (.I(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06305__A1 (.I(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06159__A1 (.I(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06877__S0 (.I(_01773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06534__S0 (.I(_01773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06419__S0 (.I(_01773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06304__S0 (.I(_01773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06158__S0 (.I(_01773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06877__S1 (.I(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06789__S1 (.I(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06701__S1 (.I(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06304__S1 (.I(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06158__S1 (.I(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06159__A2 (.I(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06393__I (.I(_01777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06313__I (.I(_01777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06185__I (.I(_01777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06174__I (.I(_01777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06161__I (.I(_01777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06899__A1 (.I(_01778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06811__A1 (.I(_01778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06422__A1 (.I(_01778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06308__A1 (.I(_01778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06166__A1 (.I(_01778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06898__S0 (.I(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06810__S0 (.I(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06722__S0 (.I(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06634__S0 (.I(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06164__S0 (.I(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06898__S1 (.I(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06810__S1 (.I(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06421__S1 (.I(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06307__S1 (.I(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06164__S1 (.I(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06899__B (.I(_01782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06811__B (.I(_01782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06422__B (.I(_01782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06308__B (.I(_01782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06166__B (.I(_01782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06847__C (.I(_01784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06759__C (.I(_01784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06671__C (.I(_01784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06583__C (.I(_01784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06168__C (.I(_01784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06192__A2 (.I(_01785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06837__A1 (.I(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06749__A1 (.I(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06661__A1 (.I(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06312__A1 (.I(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06173__A1 (.I(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06542__S0 (.I(_01787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06426__S0 (.I(_01787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06344__I (.I(_01787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06311__S0 (.I(_01787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06172__S0 (.I(_01787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06560__I (.I(_01788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06311__S1 (.I(_01788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06215__I (.I(_01788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06210__I (.I(_01788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06172__S1 (.I(_01788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06191__A1 (.I(_01790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06902__S0 (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06544__S0 (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06428__S0 (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06315__S0 (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06177__S0 (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06902__S1 (.I(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06814__S1 (.I(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06726__S1 (.I(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06638__S1 (.I(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06177__S1 (.I(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06179__A2 (.I(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06837__B (.I(_01795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06749__B (.I(_01795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06661__B (.I(_01795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06573__B (.I(_01795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06179__B (.I(_01795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06896__S0 (.I(_01798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06808__S0 (.I(_01798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06720__S0 (.I(_01798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06632__S0 (.I(_01798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06183__S0 (.I(_01798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06896__S1 (.I(_01799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06546__S1 (.I(_01799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06430__S1 (.I(_01799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06319__S1 (.I(_01799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06183__S1 (.I(_01799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06873__A1 (.I(_01802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06549__A1 (.I(_01802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06434__A1 (.I(_01802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06322__A1 (.I(_01802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06189__A1 (.I(_01802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06548__S1 (.I(_01803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06457__I (.I(_01803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06433__S1 (.I(_01803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06321__S1 (.I(_01803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06187__S1 (.I(_01803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06838__C (.I(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06750__C (.I(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06662__C (.I(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06323__C (.I(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06191__C (.I(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06192__A3 (.I(_01808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06642__B (.I(_01810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06552__B (.I(_01810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06438__B (.I(_01810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06325__B (.I(_01810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06194__B (.I(_01810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06850__S0 (.I(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06762__S0 (.I(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06674__S0 (.I(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06586__S0 (.I(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06196__I (.I(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06832__S0 (.I(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06744__S0 (.I(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06656__S0 (.I(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06555__I (.I(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06197__I (.I(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06832__S1 (.I(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06744__S1 (.I(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06326__I (.I(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06204__I (.I(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06199__I (.I(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06909__S1 (.I(_01816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06821__S1 (.I(_01816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06733__S1 (.I(_01816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06645__S1 (.I(_01816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06200__S1 (.I(_01816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06201__A2 (.I(_01817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07719__A1 (.I(_01820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07718__A1 (.I(_01820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06441__S0 (.I(_01820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06329__S0 (.I(_01820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06205__S0 (.I(_01820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07722__A1 (.I(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06556__S1 (.I(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06441__S1 (.I(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06329__S1 (.I(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06205__S1 (.I(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06207__A2 (.I(_01822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06646__B (.I(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06557__B (.I(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06442__B (.I(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06330__B (.I(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06207__B (.I(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06913__S0 (.I(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06558__S0 (.I(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06443__S0 (.I(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06332__S0 (.I(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06211__S0 (.I(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06647__S1 (.I(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06558__S1 (.I(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06443__S1 (.I(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06332__S1 (.I(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06211__S1 (.I(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06212__A2 (.I(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06219__B1 (.I(_01829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06910__A1 (.I(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06822__A1 (.I(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06734__A1 (.I(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06335__A1 (.I(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06217__A1 (.I(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06907__S0 (.I(_01831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06819__S0 (.I(_01831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06731__S0 (.I(_01831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06334__S0 (.I(_01831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06216__S0 (.I(_01831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06907__S1 (.I(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06819__S1 (.I(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06447__S1 (.I(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06334__S1 (.I(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06216__S1 (.I(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06217__A2 (.I(_01833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06220__A2 (.I(_01836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06654__S1 (.I(_01838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06566__S1 (.I(_01838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06452__S1 (.I(_01838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06339__S1 (.I(_01838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06223__S1 (.I(_01838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06224__A2 (.I(_01839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06656__S1 (.I(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06568__S1 (.I(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06454__S1 (.I(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06341__S1 (.I(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06226__S1 (.I(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06227__A2 (.I(_01842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06229__A2 (.I(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06231__A2 (.I(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06273__A2 (.I(_01848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06663__S0 (.I(_01849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06575__S0 (.I(_01849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06465__S0 (.I(_01849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06351__S0 (.I(_01849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06234__S0 (.I(_01849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06240__A2 (.I(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06244__A2 (.I(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06273__A3 (.I(_01861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06672__S0 (.I(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06584__S0 (.I(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06476__S0 (.I(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06362__S0 (.I(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06248__S0 (.I(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06249__A2 (.I(_01864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06259__A1 (.I(_01865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06252__A2 (.I(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06259__A2 (.I(_01868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06259__B1 (.I(_01870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06678__S0 (.I(_01871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06590__S0 (.I(_01871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06486__S0 (.I(_01871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06368__S0 (.I(_01871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06256__S0 (.I(_01871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06272__A2 (.I(_01875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06682__A1 (.I(_01876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06594__A1 (.I(_01876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06491__A1 (.I(_01876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06372__A1 (.I(_01876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06262__A1 (.I(_01876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06262__A2 (.I(_01877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06683__S1 (.I(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06595__S1 (.I(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06492__S1 (.I(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06374__S1 (.I(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06264__S1 (.I(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06265__A2 (.I(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06268__A2 (.I(_01883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06270__A2 (.I(_01885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06271__B2 (.I(_01886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06273__B (.I(_01888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06285__A1 (.I(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06694__S1 (.I(_01892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06606__S1 (.I(_01892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06506__S1 (.I(_01892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06391__S1 (.I(_01892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06277__S1 (.I(_01892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06278__A2 (.I(_01893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06285__A2 (.I(_01894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06696__S1 (.I(_01895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06608__S1 (.I(_01895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06509__S1 (.I(_01895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06394__S1 (.I(_01895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06280__S1 (.I(_01895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06281__A2 (.I(_01896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06283__A2 (.I(_01898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06700__C (.I(_01900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06612__C (.I(_01900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06514__C (.I(_01900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06398__C (.I(_01900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06285__C (.I(_01900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06298__A2 (.I(_01901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06287__A2 (.I(_01902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06703__S1 (.I(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06615__S1 (.I(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06517__S1 (.I(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06403__S1 (.I(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06290__S1 (.I(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06291__A2 (.I(_01906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06705__S1 (.I(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06617__S1 (.I(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06520__S1 (.I(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06405__S1 (.I(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06293__S1 (.I(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06294__A2 (.I(_01909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06297__B2 (.I(_01912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06298__A3 (.I(_01913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06325__A1 (.I(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06711__S1 (.I(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06623__S1 (.I(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06529__S1 (.I(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06412__S1 (.I(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06300__S1 (.I(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06310__A1 (.I(_01917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06310__A2 (.I(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06305__A2 (.I(_01920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06717__S0 (.I(_01922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06629__S0 (.I(_01922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06538__S0 (.I(_01922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06421__S0 (.I(_01922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06307__S0 (.I(_01922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06719__C (.I(_01925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06631__C (.I(_01925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06541__C (.I(_01925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06423__C (.I(_01925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06310__C (.I(_01925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06324__A2 (.I(_01926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06323__A1 (.I(_01928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06722__S1 (.I(_01930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06634__S1 (.I(_01930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06544__S1 (.I(_01930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06428__S1 (.I(_01930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06315__S1 (.I(_01930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06317__A2 (.I(_01931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06724__S0 (.I(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06636__S0 (.I(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06546__S0 (.I(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06430__S0 (.I(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06319__S0 (.I(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06320__A2 (.I(_01935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06731__S1 (.I(_01942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06643__S1 (.I(_01942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06553__S1 (.I(_01942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06439__S1 (.I(_01942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06327__S1 (.I(_01942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06328__A2 (.I(_01943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06330__A2 (.I(_01945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06333__A2 (.I(_01948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06336__B1 (.I(_01949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06335__A2 (.I(_01950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06337__A2 (.I(_01952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06340__A2 (.I(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06342__A2 (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06747__A1 (.I(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06659__A1 (.I(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06571__A1 (.I(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06459__A1 (.I(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06346__A1 (.I(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06746__S0 (.I(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06658__S0 (.I(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06570__S0 (.I(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06458__S0 (.I(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06345__S0 (.I(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06346__A2 (.I(_01960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06348__A2 (.I(_01962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06385__A2 (.I(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06751__S1 (.I(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06663__S1 (.I(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06575__S1 (.I(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06465__S1 (.I(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06351__S1 (.I(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06352__A2 (.I(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06753__S1 (.I(_01968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06665__S1 (.I(_01968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06577__S1 (.I(_01968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06468__S1 (.I(_01968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06354__S1 (.I(_01968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06358__A2 (.I(_01972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06360__A2 (.I(_01974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06385__A3 (.I(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06363__A2 (.I(_01977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06370__A1 (.I(_01978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06365__A2 (.I(_01979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06370__A2 (.I(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06370__B1 (.I(_01982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06375__A2 (.I(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06383__A2 (.I(_01990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06377__A2 (.I(_01991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06382__A2 (.I(_01995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06383__B2 (.I(_01997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06385__B (.I(_01999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06780__S0 (.I(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06692__S0 (.I(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06604__S0 (.I(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06504__S0 (.I(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06387__S0 (.I(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06398__A1 (.I(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06782__S0 (.I(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06694__S0 (.I(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06606__S0 (.I(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06506__S0 (.I(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06391__S0 (.I(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06392__A2 (.I(_02006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06785__A1 (.I(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06697__A1 (.I(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06609__A1 (.I(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06510__A1 (.I(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06395__A1 (.I(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06395__A2 (.I(_02009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06397__A2 (.I(_02011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06410__A2 (.I(_02013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06402__A2 (.I(_02016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06404__A2 (.I(_02018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06406__A2 (.I(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06409__B2 (.I(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06410__A3 (.I(_02024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06438__A1 (.I(_02025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06423__A1 (.I(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06801__S0 (.I(_02029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06713__S0 (.I(_02029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06625__S0 (.I(_02029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06531__S0 (.I(_02029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06415__S0 (.I(_02029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06423__A2 (.I(_02032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06803__S1 (.I(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06715__S1 (.I(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06627__S1 (.I(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06534__S1 (.I(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06419__S1 (.I(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06420__A2 (.I(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06437__A2 (.I(_02038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06808__S1 (.I(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06720__S1 (.I(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06632__S1 (.I(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06542__S1 (.I(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06426__S1 (.I(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06427__A2 (.I(_02041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06429__A2 (.I(_02043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06431__A2 (.I(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06814__S0 (.I(_02047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06726__S0 (.I(_02047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06638__S0 (.I(_02047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06548__S0 (.I(_02047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06433__S0 (.I(_02047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06434__A2 (.I(_02048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06816__C (.I(_02050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06728__C (.I(_02050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06640__C (.I(_02050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06550__C (.I(_02050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06436__C (.I(_02050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06437__A3 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06440__A2 (.I(_02054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06442__A2 (.I(_02056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06444__A2 (.I(_02058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06449__B1 (.I(_02059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06826__A1 (.I(_02060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06738__A1 (.I(_02060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06650__A1 (.I(_02060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06562__A1 (.I(_02060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06448__A1 (.I(_02060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06825__S0 (.I(_02061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06737__S0 (.I(_02061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06649__S0 (.I(_02061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06561__S0 (.I(_02061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06447__S0 (.I(_02061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06448__A2 (.I(_02062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06450__A2 (.I(_02064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06453__A2 (.I(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06456__A2 (.I(_02068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06463__A2 (.I(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06834__S1 (.I(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06746__S1 (.I(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06658__S1 (.I(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06570__S1 (.I(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06458__S1 (.I(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06459__A2 (.I(_02072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06836__S0 (.I(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06748__S0 (.I(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06660__S0 (.I(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06572__S0 (.I(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06461__S0 (.I(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06462__A2 (.I(_02075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06502__A2 (.I(_02077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06840__A1 (.I(_02078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06752__A1 (.I(_02078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06664__A1 (.I(_02078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06576__A1 (.I(_02078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06466__A1 (.I(_02078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06466__A2 (.I(_02079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06469__A2 (.I(_02082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06843__S0 (.I(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06755__S0 (.I(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06667__S0 (.I(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06579__S0 (.I(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06471__S0 (.I(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06474__A2 (.I(_02087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06502__A3 (.I(_02089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06477__A2 (.I(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06488__A1 (.I(_02091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06850__S1 (.I(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06762__S1 (.I(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06674__S1 (.I(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06586__S1 (.I(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06479__S1 (.I(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06488__B1 (.I(_02097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06855__A1 (.I(_02098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06767__A1 (.I(_02098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06679__A1 (.I(_02098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06591__A1 (.I(_02098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06487__A1 (.I(_02098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06854__S1 (.I(_02099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06766__S1 (.I(_02099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06678__S1 (.I(_02099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06590__S1 (.I(_02099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06486__S1 (.I(_02099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06857__S1 (.I(_02103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06769__S1 (.I(_02103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06681__S1 (.I(_02103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06593__S1 (.I(_02103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06490__S1 (.I(_02103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06494__A2 (.I(_02106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06500__A2 (.I(_02108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06861__S1 (.I(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06773__S1 (.I(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06685__S1 (.I(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06597__S1 (.I(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06496__S1 (.I(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06497__A2 (.I(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06499__A2 (.I(_02112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06500__B2 (.I(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06502__B (.I(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06869__A1 (.I(_02117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06781__A1 (.I(_02117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06693__A1 (.I(_02117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06605__A1 (.I(_02117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06505__A1 (.I(_02117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06514__A1 (.I(_02119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06507__A2 (.I(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06514__A2 (.I(_02121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06872__S0 (.I(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06784__S0 (.I(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06696__S0 (.I(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06608__S0 (.I(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06509__S0 (.I(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06510__A2 (.I(_02123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06513__A2 (.I(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06527__A2 (.I(_02128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06516__A2 (.I(_02129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06518__A2 (.I(_02131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06881__S0 (.I(_02133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06793__S0 (.I(_02133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06705__S0 (.I(_02133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06617__S0 (.I(_02133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06520__S0 (.I(_02133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06521__A2 (.I(_02134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06883__S0 (.I(_02136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06795__S0 (.I(_02136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06707__S0 (.I(_02136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06619__S0 (.I(_02136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06523__S0 (.I(_02136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06526__B2 (.I(_02138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06885__C (.I(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06797__C (.I(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06709__C (.I(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06621__C (.I(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06526__C (.I(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06527__A3 (.I(_02140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06552__A1 (.I(_02141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06887__S0 (.I(_02142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06799__S0 (.I(_02142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06711__S0 (.I(_02142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06623__S0 (.I(_02142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06529__S0 (.I(_02142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06541__A2 (.I(_02146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06892__A1 (.I(_02147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06804__A1 (.I(_02147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06716__A1 (.I(_02147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06628__A1 (.I(_02147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06535__A1 (.I(_02147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06535__A2 (.I(_02148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06894__A1 (.I(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06806__A1 (.I(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06718__A1 (.I(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06630__A1 (.I(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06540__A1 (.I(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06893__S1 (.I(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06805__S1 (.I(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06717__S1 (.I(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06629__S1 (.I(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06538__S1 (.I(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06551__A2 (.I(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06543__A2 (.I(_02156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06545__A2 (.I(_02158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06547__A2 (.I(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06549__A2 (.I(_02162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06551__A3 (.I(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06554__A2 (.I(_02167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06909__S0 (.I(_02169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06821__S0 (.I(_02169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06733__S0 (.I(_02169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06645__S0 (.I(_02169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06556__S0 (.I(_02169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06557__A2 (.I(_02170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06559__A2 (.I(_02172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06913__S1 (.I(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06825__S1 (.I(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06737__S1 (.I(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06649__S1 (.I(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06561__S1 (.I(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06562__A2 (.I(_02175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06564__A2 (.I(_02177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06565__B (.I(_02178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06567__A2 (.I(_02179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06569__A2 (.I(_02181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06571__A2 (.I(_02183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06573__A2 (.I(_02185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06603__A2 (.I(_02187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06576__A2 (.I(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06580__A2 (.I(_02192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06582__A2 (.I(_02194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06603__A3 (.I(_02196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06585__A2 (.I(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06587__A2 (.I(_02199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06592__A2 (.I(_02200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06592__B1 (.I(_02202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06596__A2 (.I(_02208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06601__A2 (.I(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06598__A2 (.I(_02210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06600__A2 (.I(_02212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06601__B2 (.I(_02213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06603__B (.I(_02215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06612__A1 (.I(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06607__A2 (.I(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06612__A2 (.I(_02220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06609__A2 (.I(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06611__A2 (.I(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06622__A2 (.I(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06614__A2 (.I(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06616__A2 (.I(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06618__A2 (.I(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06622__A3 (.I(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06642__A1 (.I(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06631__A2 (.I(_02239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06628__A2 (.I(_02240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06641__A2 (.I(_02244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06633__A2 (.I(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06635__A2 (.I(_02247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06640__B1 (.I(_02250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06639__A2 (.I(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06644__A2 (.I(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06646__A2 (.I(_02258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06648__A2 (.I(_02260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06650__A2 (.I(_02262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06652__A2 (.I(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06653__B (.I(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06655__A2 (.I(_02266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06657__A2 (.I(_02268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06659__A2 (.I(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06661__A2 (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06691__A2 (.I(_02274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06668__A2 (.I(_02279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06670__A2 (.I(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06691__A3 (.I(_02283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06673__A2 (.I(_02284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06680__A1 (.I(_02285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06680__A2 (.I(_02287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06680__B1 (.I(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06684__A2 (.I(_02295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06689__A2 (.I(_02296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06686__A2 (.I(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06688__A2 (.I(_02299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06689__B2 (.I(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06691__B (.I(_02302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06700__A1 (.I(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06695__A2 (.I(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06697__A2 (.I(_02308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06699__A2 (.I(_02310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06710__A2 (.I(_02312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06702__A2 (.I(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06704__A2 (.I(_02315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06706__A2 (.I(_02317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06710__A3 (.I(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06730__A1 (.I(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06712__A2 (.I(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06719__A2 (.I(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06716__A2 (.I(_02327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06729__A2 (.I(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06721__A2 (.I(_02332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06723__A2 (.I(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06728__B1 (.I(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06727__A2 (.I(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06734__A2 (.I(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06736__A2 (.I(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06738__A2 (.I(_02349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06740__A2 (.I(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06741__B (.I(_02352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06779__A2 (.I(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06756__A2 (.I(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06758__A2 (.I(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06779__A3 (.I(_02370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06761__A2 (.I(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06768__A1 (.I(_02372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06768__A2 (.I(_02374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06768__B1 (.I(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06772__A2 (.I(_02382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06774__A2 (.I(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06776__A2 (.I(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06777__B2 (.I(_02387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06779__B (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06788__A1 (.I(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06783__A2 (.I(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06785__A2 (.I(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06787__A2 (.I(_02397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06798__A2 (.I(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06790__A2 (.I(_02400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06792__A2 (.I(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06794__A2 (.I(_02404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06798__A3 (.I(_02408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06818__A1 (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06800__A2 (.I(_02410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06807__A2 (.I(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06804__A2 (.I(_02414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06817__A2 (.I(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06809__A2 (.I(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06816__A1 (.I(_02420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06811__A2 (.I(_02421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06816__B1 (.I(_02424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06815__A2 (.I(_02425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06822__A2 (.I(_02432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06824__A2 (.I(_02434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06826__A2 (.I(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06828__A2 (.I(_02438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06829__B (.I(_02439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06831__A2 (.I(_02440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06833__A2 (.I(_02442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06835__A2 (.I(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06837__A2 (.I(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06867__A2 (.I(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06844__A2 (.I(_02453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06846__A2 (.I(_02455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06867__A3 (.I(_02457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06849__A2 (.I(_02458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06856__A1 (.I(_02459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06856__A2 (.I(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06856__B1 (.I(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06860__A2 (.I(_02469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06862__A2 (.I(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06864__A2 (.I(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06865__B2 (.I(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06867__B (.I(_02476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06876__A1 (.I(_02479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06871__A2 (.I(_02480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06873__A2 (.I(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06875__A2 (.I(_02484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06886__A2 (.I(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06878__A2 (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06880__A2 (.I(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06882__A2 (.I(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06886__A3 (.I(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06906__A1 (.I(_02496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06895__A2 (.I(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06892__A2 (.I(_02501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06905__A2 (.I(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06897__A2 (.I(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06904__A1 (.I(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06904__B1 (.I(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06910__A2 (.I(_02519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06914__A2 (.I(_02523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06916__A2 (.I(_02525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06917__B (.I(_02526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06989__A1 (.I(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06919__I (.I(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10280__A1 (.I(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09518__A1 (.I(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07107__A1 (.I(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06965__A1 (.I(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06920__I (.I(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11086__A1 (.I(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10044__A1 (.I(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09966__A1 (.I(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09922__B (.I(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06921__I (.I(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10056__A2 (.I(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10040__A2 (.I(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09998__A1 (.I(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06944__A1 (.I(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06943__A1 (.I(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10447__A1 (.I(_02535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07128__A1 (.I(_02535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06928__A2 (.I(_02535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10361__A1 (.I(_02545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06967__A2 (.I(_02545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06937__I1 (.I(_02545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06982__A3 (.I(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06938__I (.I(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09648__B2 (.I(_02547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09201__A1 (.I(_02547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06975__A2 (.I(_02547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06974__A2 (.I(_02547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06939__A2 (.I(_02547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09200__A1 (.I(_02549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07097__A1 (.I(_02549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07093__A1 (.I(_02549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06947__A2 (.I(_02549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06941__A1 (.I(_02549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09202__A1 (.I(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06943__A2 (.I(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09205__B (.I(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07015__A1 (.I(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06980__A1 (.I(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06947__A1 (.I(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06946__A1 (.I(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09204__A2 (.I(_02556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07701__A2 (.I(_02556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07079__I (.I(_02556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07011__A1 (.I(_02556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06950__A1 (.I(_02556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09812__A1 (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09207__A1 (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06952__B (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06950__A2 (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09205__C (.I(_02559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07710__A2 (.I(_02559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06997__A1 (.I(_02559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06977__A1 (.I(_02559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06952__A1 (.I(_02559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06967__A1 (.I(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11111__A4 (.I(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09872__A1 (.I(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06959__A1 (.I(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09138__A1 (.I(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09126__A2 (.I(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09125__A2 (.I(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07082__A4 (.I(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06959__A2 (.I(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07003__A1 (.I(_02564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06962__B (.I(_02564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06957__I (.I(_02564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11086__A3 (.I(_02565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10252__B (.I(_02565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06979__A2 (.I(_02565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06966__A2 (.I(_02565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06959__A3 (.I(_02565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11112__A1 (.I(_02566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06959__A4 (.I(_02566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11117__A2 (.I(_02567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06967__B1 (.I(_02567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09121__I (.I(_02569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07699__A1 (.I(_02569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07021__A1 (.I(_02569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07020__A1 (.I(_02569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06962__A1 (.I(_02569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10358__A1 (.I(_02571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09858__A1 (.I(_02571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06964__A1 (.I(_02571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11105__A2 (.I(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11086__A2 (.I(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06965__A2 (.I(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07017__B (.I(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06968__B2 (.I(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11115__A2 (.I(_02576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11113__A1 (.I(_02576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06969__A2 (.I(_02576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07400__A1 (.I(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07307__A2 (.I(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07133__A1 (.I(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07038__C (.I(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06971__I (.I(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10361__A2 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09205__A2 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07096__A2 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07034__A2 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06980__A3 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09206__B2 (.I(_02589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06983__A2 (.I(_02589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06993__A2 (.I(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10183__I (.I(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07100__I (.I(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07026__A3 (.I(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06996__A2 (.I(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07038__A2 (.I(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06997__C (.I(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10042__A1 (.I(_02605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07712__A1 (.I(_02605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07118__C (.I(_02605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07016__A1 (.I(_02605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06999__B (.I(_02605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10360__I0 (.I(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07017__A1 (.I(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07117__I (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07095__A2 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07018__A2 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07009__I (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07008__A2 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09738__A1 (.I(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07092__A2 (.I(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07016__A2 (.I(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07015__A2 (.I(_02620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07014__B (.I(_02620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10043__A2 (.I(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07035__A2 (.I(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07023__A2 (.I(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10114__A2 (.I(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10039__A2 (.I(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10022__A1 (.I(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07021__A2 (.I(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10249__A2 (.I(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07099__A2 (.I(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07025__A1 (.I(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07026__A2 (.I(_02629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07024__B (.I(_02629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11094__A2 (.I(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09791__A1 (.I(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07118__A1 (.I(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07088__I (.I(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07029__A2 (.I(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07103__A3 (.I(_02635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07030__A2 (.I(_02635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10360__I1 (.I(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07037__A2 (.I(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07035__A3 (.I(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07040__I (.I(_02645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07072__A2 (.I(_02654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07053__A2 (.I(_02654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07074__A2 (.I(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07056__A2 (.I(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07076__A2 (.I(_02658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07059__A2 (.I(_02658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07078__A2 (.I(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07062__A2 (.I(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07078__A1 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07076__A1 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07074__A1 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07066__A2 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07064__A2 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09819__A1 (.I(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07125__B (.I(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07124__B (.I(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07123__B (.I(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07081__A1 (.I(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09195__A1 (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07087__A1 (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10443__A1 (.I(_02674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10039__A1 (.I(_02674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07713__A3 (.I(_02674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07112__I (.I(_02674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07086__A2 (.I(_02674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10249__A1 (.I(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10021__A1 (.I(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09778__A1 (.I(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07099__A1 (.I(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07085__A1 (.I(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10114__A1 (.I(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09794__A1 (.I(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09208__C (.I(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07091__A1 (.I(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07085__A2 (.I(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09965__A3 (.I(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09195__A2 (.I(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07086__A3 (.I(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07087__A2 (.I(_02678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09965__A1 (.I(_02679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09922__A1 (.I(_02679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07089__A1 (.I(_02679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10042__A2 (.I(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10021__B (.I(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09759__A1 (.I(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07095__A1 (.I(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07091__A2 (.I(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10024__A2 (.I(_02682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10023__C (.I(_02682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07097__A3 (.I(_02682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07093__A4 (.I(_02682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11098__C (.I(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11094__A1 (.I(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10112__A1 (.I(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07712__C (.I(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07096__A1 (.I(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10253__A1 (.I(_02690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10228__I (.I(_02690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10217__I (.I(_02690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10206__I (.I(_02690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07101__I (.I(_02690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10251__B2 (.I(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10248__B (.I(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10247__A2 (.I(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10246__A2 (.I(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07102__B (.I(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11122__A1 (.I(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11106__A1 (.I(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11098__B (.I(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11089__A1 (.I(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07105__A1 (.I(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07699__A2 (.I(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07119__I (.I(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07107__A2 (.I(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10283__A2 (.I(_02696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07111__B (.I(_02696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07108__B (.I(_02696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10182__A1 (.I(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10181__A2 (.I(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09140__B (.I(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07121__B (.I(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07113__A2 (.I(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10468__A1 (.I(_02700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10455__I1 (.I(_02700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10365__A1 (.I(_02700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07429__A1 (.I(_02700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07116__A2 (.I(_02700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10473__A1 (.I(_02701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10464__A1 (.I(_02701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07215__A1 (.I(_02701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07148__A1 (.I(_02701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07116__A3 (.I(_02701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10021__A2 (.I(_02703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09965__A2 (.I(_02703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09922__A2 (.I(_02703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09208__A1 (.I(_02703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07118__A2 (.I(_02703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10443__A2 (.I(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07120__B (.I(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10280__A2 (.I(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10256__A2 (.I(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10248__A2 (.I(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10122__A2 (.I(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07120__C (.I(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07209__A1 (.I(_02708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07129__A1 (.I(_02708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07209__A2 (.I(_02710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07129__A2 (.I(_02710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07400__A2 (.I(_02714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07133__A2 (.I(_02714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07524__A1 (.I(_02716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07364__A1 (.I(_02716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07237__A1 (.I(_02716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07140__A1 (.I(_02716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07341__A1 (.I(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07279__A2 (.I(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07138__I (.I(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11230__A1 (.I(_02722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09873__A1 (.I(_02722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09255__A1 (.I(_02722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08857__A1 (.I(_02722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07141__I (.I(_02722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10405__A1 (.I(_02723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08010__A1 (.I(_02723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07651__A1 (.I(_02723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07259__A1 (.I(_02723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07150__A1 (.I(_02723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07816__A1 (.I(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07525__A3 (.I(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07305__A2 (.I(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07147__A2 (.I(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07143__A2 (.I(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07307__A1 (.I(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07200__A1 (.I(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07168__I (.I(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07154__I (.I(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07145__A1 (.I(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11270__A1 (.I(_02730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10898__I (.I(_02730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09214__I (.I(_02730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07149__I (.I(_02730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09168__A1 (.I(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09147__A1 (.I(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07366__A1 (.I(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07239__A1 (.I(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07150__A2 (.I(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07204__A2 (.I(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07173__I (.I(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07159__I (.I(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07151__I (.I(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07187__A1 (.I(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07181__A1 (.I(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07175__A1 (.I(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07167__A1 (.I(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07161__A1 (.I(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07337__S (.I(_02734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07201__A1 (.I(_02734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07195__A1 (.I(_02734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07189__A1 (.I(_02734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07153__I (.I(_02734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07333__S (.I(_02736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07329__S (.I(_02736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07302__I (.I(_02736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07162__A1 (.I(_02736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07155__A2 (.I(_02736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10125__I (.I(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08916__I (.I(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08267__I (.I(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07157__I (.I(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11124__I (.I(_02739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10977__I (.I(_02739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07613__I (.I(_02739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07362__I (.I(_02739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07158__I (.I(_02739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07286__A1 (.I(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07263__A1 (.I(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07243__A1 (.I(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07221__A1 (.I(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07161__A2 (.I(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07205__A1 (.I(_02741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07199__A1 (.I(_02741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07193__A1 (.I(_02741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07166__A2 (.I(_02741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07160__A2 (.I(_02741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10132__I (.I(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08923__I (.I(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08274__I (.I(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07164__I (.I(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11130__I (.I(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10983__I (.I(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07622__I (.I(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07371__I (.I(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07165__I (.I(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07288__A1 (.I(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07265__A1 (.I(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07245__A1 (.I(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07223__A1 (.I(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07167__A2 (.I(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07194__A1 (.I(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07188__A1 (.I(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07182__A1 (.I(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07176__A1 (.I(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07169__A1 (.I(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10136__I (.I(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08927__I (.I(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08278__I (.I(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07171__I (.I(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11133__I (.I(_02751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10986__I (.I(_02751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07626__I (.I(_02751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07375__I (.I(_02751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07172__I (.I(_02751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07291__A1 (.I(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07268__A1 (.I(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07248__A1 (.I(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07226__A1 (.I(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07175__A2 (.I(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07198__A2 (.I(_02753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07192__A2 (.I(_02753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07186__A2 (.I(_02753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07180__A2 (.I(_02753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07174__A2 (.I(_02753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10141__I (.I(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08932__I (.I(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08283__I (.I(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07178__I (.I(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11137__I (.I(_02757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10990__I (.I(_02757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07631__I (.I(_02757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07380__I (.I(_02757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07179__I (.I(_02757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07293__A1 (.I(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07270__A1 (.I(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07250__A1 (.I(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07228__A1 (.I(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07181__A2 (.I(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10145__I (.I(_02761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08936__I (.I(_02761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08287__I (.I(_02761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07184__I (.I(_02761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11140__I (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10993__I (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07635__I (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07384__I (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07185__I (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07295__A1 (.I(_02763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07272__A1 (.I(_02763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07252__A1 (.I(_02763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07230__A1 (.I(_02763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07187__A2 (.I(_02763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10149__I (.I(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08940__I (.I(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08291__I (.I(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07190__I (.I(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11143__I (.I(_02767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10996__I (.I(_02767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07639__I (.I(_02767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07388__I (.I(_02767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07191__I (.I(_02767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07297__A1 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07274__A1 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07254__A1 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07232__A1 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07193__A2 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10153__I (.I(_02771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08944__I (.I(_02771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08295__I (.I(_02771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07196__I (.I(_02771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11146__I (.I(_02772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10999__I (.I(_02772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07643__I (.I(_02772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07392__I (.I(_02772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07197__I (.I(_02772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07299__A1 (.I(_02773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07276__A1 (.I(_02773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07256__A1 (.I(_02773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07234__A1 (.I(_02773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07199__A2 (.I(_02773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10157__I (.I(_02776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08948__I (.I(_02776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08299__I (.I(_02776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07202__I (.I(_02776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11149__I (.I(_02777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11002__I (.I(_02777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07647__I (.I(_02777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07396__I (.I(_02777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07203__I (.I(_02777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07301__A1 (.I(_02778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07278__A1 (.I(_02778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07258__A1 (.I(_02778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07236__A1 (.I(_02778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07205__A2 (.I(_02778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07949__A2 (.I(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07342__A1 (.I(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07280__A1 (.I(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07211__A2 (.I(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10878__A1 (.I(_02785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10633__A1 (.I(_02785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09275__A1 (.I(_02785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09081__A1 (.I(_02785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07212__I (.I(_02785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10957__A2 (.I(_02786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08790__A1 (.I(_02786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08343__A1 (.I(_02786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08209__A1 (.I(_02786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07217__A1 (.I(_02786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11290__A1 (.I(_02789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10576__I (.I(_02789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08078__I (.I(_02789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07216__I (.I(_02789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07235__A2 (.I(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07224__I (.I(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07219__I (.I(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07218__I (.I(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07230__A2 (.I(_02792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07228__A2 (.I(_02792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07226__A2 (.I(_02792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07223__A2 (.I(_02792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07221__A2 (.I(_02792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07233__A2 (.I(_02796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07231__A2 (.I(_02796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07229__A2 (.I(_02796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07227__A2 (.I(_02796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07225__A2 (.I(_02796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10484__A1 (.I(_02803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09650__A1 (.I(_02803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09496__A1 (.I(_02803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08708__A1 (.I(_02803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07238__I (.I(_02803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08031__A1 (.I(_02804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07818__A1 (.I(_02804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07744__A2 (.I(_02804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07309__A1 (.I(_02804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07239__A2 (.I(_02804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07257__A2 (.I(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07246__I (.I(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07241__I (.I(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07240__I (.I(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07252__A2 (.I(_02806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07250__A2 (.I(_02806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07248__A2 (.I(_02806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07245__A2 (.I(_02806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07243__A2 (.I(_02806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07258__A2 (.I(_02807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07256__A2 (.I(_02807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07254__A2 (.I(_02807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07244__A2 (.I(_02807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07242__A2 (.I(_02807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07255__A2 (.I(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07253__A2 (.I(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07251__A2 (.I(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07249__A2 (.I(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07247__A2 (.I(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07277__A2 (.I(_02817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07266__I (.I(_02817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07261__I (.I(_02817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07260__I (.I(_02817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07272__A2 (.I(_02818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07270__A2 (.I(_02818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07268__A2 (.I(_02818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07265__A2 (.I(_02818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07263__A2 (.I(_02818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07278__A2 (.I(_02819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07276__A2 (.I(_02819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07274__A2 (.I(_02819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07264__A2 (.I(_02819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07262__A2 (.I(_02819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07275__A2 (.I(_02822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07273__A2 (.I(_02822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07271__A2 (.I(_02822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07269__A2 (.I(_02822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07267__A2 (.I(_02822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11250__A1 (.I(_02830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09476__A1 (.I(_02830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09101__A1 (.I(_02830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08817__A1 (.I(_02830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07281__I (.I(_02830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10899__A2 (.I(_02831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08363__A1 (.I(_02831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07969__A1 (.I(_02831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07671__A1 (.I(_02831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07282__A2 (.I(_02831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07300__A2 (.I(_02832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07289__I (.I(_02832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07284__I (.I(_02832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07283__I (.I(_02832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07295__A2 (.I(_02833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07293__A2 (.I(_02833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07291__A2 (.I(_02833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07288__A2 (.I(_02833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07286__A2 (.I(_02833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07298__A2 (.I(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07296__A2 (.I(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07294__A2 (.I(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07292__A2 (.I(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07290__A2 (.I(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07325__S (.I(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07321__S (.I(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07317__S (.I(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07313__S (.I(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07303__S (.I(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11214__I0 (.I(_02845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09363__I (.I(_02845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08383__I (.I(_02845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07304__I (.I(_02845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11212__A1 (.I(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08877__I (.I(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07948__I (.I(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07308__I (.I(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10405__A2 (.I(_02850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08209__A2 (.I(_02850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07671__A2 (.I(_02850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07344__A1 (.I(_02850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07309__A2 (.I(_02850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07339__S (.I(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07335__S (.I(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07331__S (.I(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07310__I (.I(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07327__S (.I(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07323__S (.I(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07319__S (.I(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07315__S (.I(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07311__S (.I(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11216__I0 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09368__I (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08388__I (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07314__I (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08213__I0 (.I(_02855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07955__I0 (.I(_02855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07675__I0 (.I(_02855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07348__I0 (.I(_02855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07315__I0 (.I(_02855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11218__I0 (.I(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09371__I (.I(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08391__I (.I(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07318__I (.I(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08215__I0 (.I(_02858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07957__I0 (.I(_02858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07677__I0 (.I(_02858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07350__I0 (.I(_02858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07319__I0 (.I(_02858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11220__I0 (.I(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09374__I (.I(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08394__I (.I(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07322__I (.I(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08217__I0 (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07959__I0 (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07679__I0 (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07352__I0 (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07323__I0 (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11222__I0 (.I(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09377__I (.I(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08397__I (.I(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07326__I (.I(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08219__I0 (.I(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07961__I0 (.I(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07681__I0 (.I(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07354__I0 (.I(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07327__I0 (.I(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11224__I0 (.I(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09380__I (.I(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08400__I (.I(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07330__I (.I(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08221__I0 (.I(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07963__I0 (.I(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07683__I0 (.I(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07356__I0 (.I(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07331__I0 (.I(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11226__I0 (.I(_02869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09383__I (.I(_02869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08403__I (.I(_02869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07334__I (.I(_02869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08223__I0 (.I(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07965__I0 (.I(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07685__I0 (.I(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07358__I0 (.I(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07335__I0 (.I(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11228__I0 (.I(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09386__I (.I(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08406__I (.I(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07338__I (.I(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08225__I0 (.I(_02873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07967__I0 (.I(_02873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07687__I0 (.I(_02873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07360__I0 (.I(_02873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07339__I0 (.I(_02873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10681__A1 (.I(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08748__A1 (.I(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08660__A1 (.I(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08554__A1 (.I(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07343__I (.I(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11290__A2 (.I(_02877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11045__A2 (.I(_02877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08303__A1 (.I(_02877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07789__A1 (.I(_02877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07344__A2 (.I(_02877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07360__S (.I(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07358__S (.I(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07356__S (.I(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07345__I (.I(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07354__S (.I(_02879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07352__S (.I(_02879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07350__S (.I(_02879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07348__S (.I(_02879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07346__S (.I(_02879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11294__A1 (.I(_02888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11274__A1 (.I(_02888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11254__A1 (.I(_02888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07494__I (.I(_02888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07363__I (.I(_02888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07478__A1 (.I(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07455__A1 (.I(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07435__A1 (.I(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07410__A1 (.I(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07370__A1 (.I(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10551__A1 (.I(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10127__A1 (.I(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09407__A1 (.I(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08918__A1 (.I(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07365__I (.I(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11212__A2 (.I(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08058__A1 (.I(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07724__A2 (.I(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07593__A1 (.I(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07366__A2 (.I(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07387__A2 (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07383__A2 (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07379__A2 (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07374__A2 (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07370__A2 (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07399__A2 (.I(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07395__A2 (.I(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07391__A2 (.I(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07373__A2 (.I(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07369__A2 (.I(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11296__A1 (.I(_02896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11276__A1 (.I(_02896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11256__A1 (.I(_02896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07502__I (.I(_02896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07372__I (.I(_02896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07480__A1 (.I(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07457__A1 (.I(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07437__A1 (.I(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07412__A1 (.I(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07374__A1 (.I(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11299__A1 (.I(_02899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11279__A1 (.I(_02899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11259__A1 (.I(_02899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07505__I (.I(_02899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07376__I (.I(_02899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07483__A1 (.I(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07460__A1 (.I(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07440__A1 (.I(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07415__A1 (.I(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07379__A1 (.I(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07394__A2 (.I(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07390__A2 (.I(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07386__A2 (.I(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07382__A2 (.I(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07378__A2 (.I(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11301__A1 (.I(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11281__A1 (.I(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11261__A1 (.I(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07509__I (.I(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07381__I (.I(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07485__A1 (.I(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07462__A1 (.I(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07442__A1 (.I(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07417__A1 (.I(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07383__A1 (.I(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11303__A1 (.I(_02906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11283__A1 (.I(_02906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11263__A1 (.I(_02906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07512__I (.I(_02906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07385__I (.I(_02906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07487__A1 (.I(_02907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07464__A1 (.I(_02907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07444__A1 (.I(_02907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07419__A1 (.I(_02907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07387__A1 (.I(_02907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11305__A1 (.I(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11285__A1 (.I(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11265__A1 (.I(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07515__I (.I(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07389__I (.I(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07489__A1 (.I(_02910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07466__A1 (.I(_02910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07446__A1 (.I(_02910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07421__A1 (.I(_02910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07391__A1 (.I(_02910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11307__A1 (.I(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11287__A1 (.I(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11267__A1 (.I(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07518__I (.I(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07393__I (.I(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07491__A1 (.I(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07468__A1 (.I(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07448__A1 (.I(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07423__A1 (.I(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07395__A1 (.I(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11309__A1 (.I(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11289__A1 (.I(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11269__A1 (.I(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07521__I (.I(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07397__I (.I(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07493__A1 (.I(_02916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07470__A1 (.I(_02916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07450__A1 (.I(_02916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07425__A1 (.I(_02916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07399__A1 (.I(_02916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07615__A2 (.I(_02919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07495__A2 (.I(_02919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07472__A2 (.I(_02919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07402__A2 (.I(_02919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10978__A1 (.I(_02920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08972__A1 (.I(_02920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08428__A1 (.I(_02920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08120__A1 (.I(_02920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07403__I (.I(_02920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10511__A2 (.I(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10260__A2 (.I(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08622__A2 (.I(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07451__A1 (.I(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07406__A1 (.I(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10742__A1 (.I(_02922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07927__I (.I(_02922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07858__I (.I(_02922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07405__I (.I(_02922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08058__A2 (.I(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08031__A2 (.I(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08010__A2 (.I(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07969__A2 (.I(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07406__A2 (.I(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07419__A2 (.I(_02925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07417__A2 (.I(_02925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07415__A2 (.I(_02925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07412__A2 (.I(_02925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07410__A2 (.I(_02925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07425__A2 (.I(_02926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07423__A2 (.I(_02926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07421__A2 (.I(_02926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07411__A2 (.I(_02926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07409__A2 (.I(_02926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07422__A2 (.I(_02929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07420__A2 (.I(_02929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07418__A2 (.I(_02929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07416__A2 (.I(_02929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07414__A2 (.I(_02929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07764__A2 (.I(_02936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07571__A2 (.I(_02936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07549__A2 (.I(_02936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07427__A2 (.I(_02936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10789__A1 (.I(_02937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09428__A1 (.I(_02937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08640__A1 (.I(_02937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08227__A1 (.I(_02937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07428__I (.I(_02937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11152__A2 (.I(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10939__A2 (.I(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09168__A2 (.I(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07879__A2 (.I(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07431__A1 (.I(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09235__A1 (.I(_02939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07548__I (.I(_02939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07471__I (.I(_02939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07430__I (.I(_02939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09101__A2 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09081__A2 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08660__A2 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07451__A2 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07431__A2 (.I(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07444__A2 (.I(_02942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07442__A2 (.I(_02942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07440__A2 (.I(_02942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07437__A2 (.I(_02942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07435__A2 (.I(_02942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07447__A2 (.I(_02946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07445__A2 (.I(_02946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07443__A2 (.I(_02946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07441__A2 (.I(_02946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07439__A2 (.I(_02946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07464__A2 (.I(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07462__A2 (.I(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07460__A2 (.I(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07457__A2 (.I(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07455__A2 (.I(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10127__A2 (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09496__A2 (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09255__A2 (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07497__A1 (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07474__A1 (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10367__A1 (.I(_02966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08992__A1 (.I(_02966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08455__A1 (.I(_02966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08141__A1 (.I(_02966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07473__I (.I(_02966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10423__A2 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08495__A2 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08079__A2 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07859__A2 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07474__A2 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07487__A2 (.I(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07485__A2 (.I(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07483__A2 (.I(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07480__A2 (.I(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07478__A2 (.I(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07493__A2 (.I(_02970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07491__A2 (.I(_02970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07489__A2 (.I(_02970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07479__A2 (.I(_02970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07477__A2 (.I(_02970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07490__A2 (.I(_02973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07488__A2 (.I(_02973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07486__A2 (.I(_02973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07484__A2 (.I(_02973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07482__A2 (.I(_02973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07597__A1 (.I(_02980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07577__A1 (.I(_02980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07555__A1 (.I(_02980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07532__A1 (.I(_02980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07501__A1 (.I(_02980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10851__A1 (.I(_02981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09012__A1 (.I(_02981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08475__A1 (.I(_02981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08169__A1 (.I(_02981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07496__I (.I(_02981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10577__A2 (.I(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09215__A2 (.I(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08878__A2 (.I(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07900__A2 (.I(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07497__A2 (.I(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07514__A2 (.I(_02984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07511__A2 (.I(_02984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07508__A2 (.I(_02984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07504__A2 (.I(_02984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07501__A2 (.I(_02984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07523__A2 (.I(_02985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07520__A2 (.I(_02985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07517__A2 (.I(_02985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07503__A2 (.I(_02985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07500__A2 (.I(_02985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07599__A1 (.I(_02987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07579__A1 (.I(_02987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07557__A1 (.I(_02987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07534__A1 (.I(_02987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07504__A1 (.I(_02987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07602__A1 (.I(_02989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07582__A1 (.I(_02989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07560__A1 (.I(_02989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07537__A1 (.I(_02989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07508__A1 (.I(_02989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07519__A2 (.I(_02990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07516__A2 (.I(_02990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07513__A2 (.I(_02990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07510__A2 (.I(_02990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07507__A2 (.I(_02990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07604__A1 (.I(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07584__A1 (.I(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07562__A1 (.I(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07539__A1 (.I(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07511__A1 (.I(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07606__A1 (.I(_02994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07586__A1 (.I(_02994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07564__A1 (.I(_02994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07541__A1 (.I(_02994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07514__A1 (.I(_02994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07608__A1 (.I(_02996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07588__A1 (.I(_02996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07566__A1 (.I(_02996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07543__A1 (.I(_02996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07517__A1 (.I(_02996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07610__A1 (.I(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07590__A1 (.I(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07568__A1 (.I(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07545__A1 (.I(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07520__A1 (.I(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07612__A1 (.I(_03000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07592__A1 (.I(_03000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07570__A1 (.I(_03000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07547__A1 (.I(_03000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07523__A1 (.I(_03000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10721__A1 (.I(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09449__A1 (.I(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08837__A1 (.I(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07989__I (.I(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07528__A1 (.I(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10919__A1 (.I(_03004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08168__I (.I(_03004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08099__I (.I(_03004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07527__I (.I(_03004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08141__A2 (.I(_03005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08120__A2 (.I(_03005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07651__A2 (.I(_03005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07593__A2 (.I(_03005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07528__A2 (.I(_03005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07546__A2 (.I(_03006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07535__I (.I(_03006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07530__I (.I(_03006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07529__I (.I(_03006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07541__A2 (.I(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07539__A2 (.I(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07537__A2 (.I(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07534__A2 (.I(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07532__A2 (.I(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07547__A2 (.I(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07545__A2 (.I(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07543__A2 (.I(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07533__A2 (.I(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07531__A2 (.I(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07544__A2 (.I(_03011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07542__A2 (.I(_03011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07540__A2 (.I(_03011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07538__A2 (.I(_03011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07536__A2 (.I(_03011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09061__A1 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07766__A1 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07617__A1 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07573__A1 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07551__A1 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11270__A2 (.I(_03019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10769__A1 (.I(_03019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09343__A1 (.I(_03019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08681__A1 (.I(_03019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07550__I (.I(_03019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11172__A2 (.I(_03020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08533__A2 (.I(_03020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08384__A2 (.I(_03020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08247__A2 (.I(_03020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07551__A2 (.I(_03020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11125__A2 (.I(_03033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10810__A1 (.I(_03033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09034__A1 (.I(_03033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07838__A1 (.I(_03033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07572__I (.I(_03033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10919__A2 (.I(_03034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09389__A2 (.I(_03034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09147__A2 (.I(_03034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07928__A2 (.I(_03034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07573__A2 (.I(_03034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07586__A2 (.I(_03036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07584__A2 (.I(_03036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07582__A2 (.I(_03036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07579__A2 (.I(_03036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07577__A2 (.I(_03036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07592__A2 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07590__A2 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07588__A2 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07578__A2 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07576__A2 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07589__A2 (.I(_03040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07587__A2 (.I(_03040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07585__A2 (.I(_03040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07583__A2 (.I(_03040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07581__A2 (.I(_03040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07611__A2 (.I(_03047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07600__I (.I(_03047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07595__I (.I(_03047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07594__I (.I(_03047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07606__A2 (.I(_03048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07604__A2 (.I(_03048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07602__A2 (.I(_03048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07599__A2 (.I(_03048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07597__A2 (.I(_03048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07612__A2 (.I(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07610__A2 (.I(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07608__A2 (.I(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07598__A2 (.I(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07596__A2 (.I(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07609__A2 (.I(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07607__A2 (.I(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07605__A2 (.I(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07603__A2 (.I(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07601__A2 (.I(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08140__I (.I(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08030__I (.I(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07899__I (.I(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07786__I (.I(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07614__I (.I(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07770__A1 (.I(_03060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07748__A1 (.I(_03060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07728__A1 (.I(_03060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07655__A1 (.I(_03060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07621__A1 (.I(_03060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11025__A1 (.I(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10742__A2 (.I(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08952__A1 (.I(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08602__A1 (.I(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07616__I (.I(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10531__A2 (.I(_03062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10161__A2 (.I(_03062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08409__A2 (.I(_03062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08100__A2 (.I(_03062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07617__A2 (.I(_03062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07638__A2 (.I(_03064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07634__A2 (.I(_03064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07630__A2 (.I(_03064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07625__A2 (.I(_03064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07621__A2 (.I(_03064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08146__I (.I(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08036__I (.I(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07905__I (.I(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07794__I (.I(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07623__I (.I(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07772__A1 (.I(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07750__A1 (.I(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07730__A1 (.I(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07657__A1 (.I(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07625__A1 (.I(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08149__I (.I(_03070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08039__I (.I(_03070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07908__I (.I(_03070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07797__I (.I(_03070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07627__I (.I(_03070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07775__A1 (.I(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07753__A1 (.I(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07733__A1 (.I(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07660__A1 (.I(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07630__A1 (.I(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07645__A2 (.I(_03072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07641__A2 (.I(_03072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07637__A2 (.I(_03072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07633__A2 (.I(_03072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07629__A2 (.I(_03072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08153__I (.I(_03074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08043__I (.I(_03074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07912__I (.I(_03074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07801__I (.I(_03074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07632__I (.I(_03074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07777__A1 (.I(_03075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07755__A1 (.I(_03075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07735__A1 (.I(_03075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07662__A1 (.I(_03075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07634__A1 (.I(_03075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08156__I (.I(_03077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08046__I (.I(_03077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07915__I (.I(_03077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07804__I (.I(_03077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07636__I (.I(_03077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07779__A1 (.I(_03078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07757__A1 (.I(_03078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07737__A1 (.I(_03078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07664__A1 (.I(_03078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07638__A1 (.I(_03078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08159__I (.I(_03080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08049__I (.I(_03080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07918__I (.I(_03080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07807__I (.I(_03080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07640__I (.I(_03080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07781__A1 (.I(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07759__A1 (.I(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07739__A1 (.I(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07666__A1 (.I(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07642__A1 (.I(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08162__I (.I(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08052__I (.I(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07921__I (.I(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07810__I (.I(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07644__I (.I(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07783__A1 (.I(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07761__A1 (.I(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07741__A1 (.I(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07668__A1 (.I(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07646__A1 (.I(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08165__I (.I(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08055__I (.I(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07924__I (.I(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07813__I (.I(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07648__I (.I(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07785__A1 (.I(_03087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07763__A1 (.I(_03087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07743__A1 (.I(_03087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07670__A1 (.I(_03087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07650__A1 (.I(_03087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07669__A2 (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07658__I (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07653__I (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07652__I (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07664__A2 (.I(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07662__A2 (.I(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07660__A2 (.I(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07657__A2 (.I(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07655__A2 (.I(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07687__S (.I(_03101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07685__S (.I(_03101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07683__S (.I(_03101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07672__I (.I(_03101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07681__S (.I(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07679__S (.I(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07677__S (.I(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07675__S (.I(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07673__S (.I(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11123__A1 (.I(_03111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09197__A1 (.I(_03111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09127__A1 (.I(_03111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09123__A1 (.I(_03111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07690__I (.I(_03111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10575__A1 (.I(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09213__A1 (.I(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09144__A1 (.I(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09135__A1 (.I(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07698__A1 (.I(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09706__A1 (.I(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09698__A1 (.I(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09690__A1 (.I(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09679__I (.I(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07693__I (.I(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10002__A1 (.I(_03115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09995__A1 (.I(_03115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09990__A1 (.I(_03115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09968__A1 (.I(_03115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07695__A1 (.I(_03115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10630__S (.I(_03116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10619__I (.I(_03116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10608__I (.I(_03116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10597__I (.I(_03116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07695__B (.I(_03116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10444__A1 (.I(_03118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09838__A1 (.I(_03118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09796__I (.I(_03118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09771__A1 (.I(_03118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07697__B (.I(_03118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11320__A1 (.I(_03119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07720__A1 (.I(_03119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07714__A1 (.I(_03119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07698__A2 (.I(_03119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10253__A2 (.I(_03123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10252__C (.I(_03123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10250__A2 (.I(_03123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09122__A2 (.I(_03123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07703__A2 (.I(_03123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09557__A1 (.I(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09536__I (.I(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09525__I (.I(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07712__B (.I(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07737__A2 (.I(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07735__A2 (.I(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07733__A2 (.I(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07730__A2 (.I(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07728__A2 (.I(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07743__A2 (.I(_03143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07741__A2 (.I(_03143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07739__A2 (.I(_03143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07729__A2 (.I(_03143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07727__A2 (.I(_03143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07740__A2 (.I(_03146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07738__A2 (.I(_03146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07736__A2 (.I(_03146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07734__A2 (.I(_03146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07732__A2 (.I(_03146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07757__A2 (.I(_03154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07755__A2 (.I(_03154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07753__A2 (.I(_03154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07750__A2 (.I(_03154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07748__A2 (.I(_03154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07763__A2 (.I(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07761__A2 (.I(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07759__A2 (.I(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07749__A2 (.I(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07747__A2 (.I(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07760__A2 (.I(_03158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07758__A2 (.I(_03158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07756__A2 (.I(_03158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07754__A2 (.I(_03158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07752__A2 (.I(_03158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11192__A2 (.I(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10701__A1 (.I(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09296__A1 (.I(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08728__A1 (.I(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07765__I (.I(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11065__A2 (.I(_03166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09364__A2 (.I(_03166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08513__A2 (.I(_03166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08269__A2 (.I(_03166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07766__A2 (.I(_03166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07779__A2 (.I(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07777__A2 (.I(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07775__A2 (.I(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07772__A2 (.I(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07770__A2 (.I(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07782__A2 (.I(_03172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07780__A2 (.I(_03172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07778__A2 (.I(_03172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07776__A2 (.I(_03172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07774__A2 (.I(_03172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07883__A1 (.I(_03179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07863__A1 (.I(_03179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07842__A1 (.I(_03179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07822__A1 (.I(_03179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07793__A1 (.I(_03179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09427__I (.I(_03180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09323__A1 (.I(_03180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09033__I (.I(_03180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07788__I (.I(_03180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09012__A2 (.I(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08992__A2 (.I(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08972__A2 (.I(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08952__A2 (.I(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07789__A2 (.I(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07885__A1 (.I(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07865__A1 (.I(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07844__A1 (.I(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07824__A1 (.I(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07796__A1 (.I(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07888__A1 (.I(_03188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07868__A1 (.I(_03188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07847__A1 (.I(_03188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07827__A1 (.I(_03188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07800__A1 (.I(_03188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07890__A1 (.I(_03191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07870__A1 (.I(_03191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07849__A1 (.I(_03191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07829__A1 (.I(_03191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07803__A1 (.I(_03191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07892__A1 (.I(_03193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07872__A1 (.I(_03193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07851__A1 (.I(_03193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07831__A1 (.I(_03193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07806__A1 (.I(_03193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07894__A1 (.I(_03195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07874__A1 (.I(_03195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07853__A1 (.I(_03195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07833__A1 (.I(_03195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07809__A1 (.I(_03195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07896__A1 (.I(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07876__A1 (.I(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07855__A1 (.I(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07835__A1 (.I(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07812__A1 (.I(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07898__A1 (.I(_03199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07878__A1 (.I(_03199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07857__A1 (.I(_03199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07837__A1 (.I(_03199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07815__A1 (.I(_03199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08789__I (.I(_03201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08768__A1 (.I(_03201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08601__I (.I(_03201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07817__I (.I(_03201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08475__A2 (.I(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08455__A2 (.I(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08428__A2 (.I(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07838__A2 (.I(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07818__A2 (.I(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07837__A2 (.I(_03205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07835__A2 (.I(_03205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07833__A2 (.I(_03205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07823__A2 (.I(_03205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07821__A2 (.I(_03205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07834__A2 (.I(_03208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07832__A2 (.I(_03208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07830__A2 (.I(_03208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07828__A2 (.I(_03208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07826__A2 (.I(_03208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07856__A2 (.I(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07845__I (.I(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07840__I (.I(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07839__I (.I(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07857__A2 (.I(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07855__A2 (.I(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07853__A2 (.I(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07843__A2 (.I(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07841__A2 (.I(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07854__A2 (.I(_03220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07852__A2 (.I(_03220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07850__A2 (.I(_03220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07848__A2 (.I(_03220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07846__A2 (.I(_03220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10878__A2 (.I(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08554__A2 (.I(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07900__A1 (.I(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07879__A1 (.I(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07859__A1 (.I(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07877__A2 (.I(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07866__I (.I(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07861__I (.I(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07860__I (.I(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07872__A2 (.I(_03229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07870__A2 (.I(_03229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07868__A2 (.I(_03229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07865__A2 (.I(_03229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07863__A2 (.I(_03229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07878__A2 (.I(_03230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07876__A2 (.I(_03230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07874__A2 (.I(_03230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07864__A2 (.I(_03230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07862__A2 (.I(_03230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07875__A2 (.I(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07873__A2 (.I(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07871__A2 (.I(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07869__A2 (.I(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07867__A2 (.I(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07892__A2 (.I(_03241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07890__A2 (.I(_03241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07888__A2 (.I(_03241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07885__A2 (.I(_03241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07883__A2 (.I(_03241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07898__A2 (.I(_03242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07896__A2 (.I(_03242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07894__A2 (.I(_03242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07884__A2 (.I(_03242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07882__A2 (.I(_03242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07895__A2 (.I(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07893__A2 (.I(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07891__A2 (.I(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07889__A2 (.I(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07887__A2 (.I(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08014__A1 (.I(_03252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07994__A1 (.I(_03252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07973__A1 (.I(_03252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07932__A1 (.I(_03252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07904__A1 (.I(_03252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07925__A2 (.I(_03253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07909__I (.I(_03253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07902__I (.I(_03253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07901__I (.I(_03253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07917__A2 (.I(_03254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07914__A2 (.I(_03254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07911__A2 (.I(_03254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07907__A2 (.I(_03254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07904__A2 (.I(_03254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07926__A2 (.I(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07923__A2 (.I(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07920__A2 (.I(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07906__A2 (.I(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07903__A2 (.I(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08016__A1 (.I(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07996__A1 (.I(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07975__A1 (.I(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07934__A1 (.I(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07907__A1 (.I(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08019__A1 (.I(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07999__A1 (.I(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07978__A1 (.I(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07937__A1 (.I(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07911__A1 (.I(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07922__A2 (.I(_03260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07919__A2 (.I(_03260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07916__A2 (.I(_03260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07913__A2 (.I(_03260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07910__A2 (.I(_03260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08021__A1 (.I(_03262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08001__A1 (.I(_03262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07980__A1 (.I(_03262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07939__A1 (.I(_03262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07914__A1 (.I(_03262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08023__A1 (.I(_03264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08003__A1 (.I(_03264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07982__A1 (.I(_03264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07941__A1 (.I(_03264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07917__A1 (.I(_03264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08025__A1 (.I(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08005__A1 (.I(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07984__A1 (.I(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07943__A1 (.I(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07920__A1 (.I(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08027__A1 (.I(_03268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08007__A1 (.I(_03268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07986__A1 (.I(_03268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07945__A1 (.I(_03268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07923__A1 (.I(_03268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08029__A1 (.I(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08009__A1 (.I(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07988__A1 (.I(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07947__A1 (.I(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07926__A1 (.I(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08581__A1 (.I(_03272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08533__A1 (.I(_03272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08513__A1 (.I(_03272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07990__A1 (.I(_03272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07928__A1 (.I(_03272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07941__A2 (.I(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07939__A2 (.I(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07937__A2 (.I(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07934__A2 (.I(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07932__A2 (.I(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07947__A2 (.I(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07945__A2 (.I(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07943__A2 (.I(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07933__A2 (.I(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07931__A2 (.I(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07944__A2 (.I(_03278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07942__A2 (.I(_03278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07940__A2 (.I(_03278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07938__A2 (.I(_03278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07936__A2 (.I(_03278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08622__A1 (.I(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08495__A1 (.I(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08409__A1 (.I(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08384__A1 (.I(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07951__A1 (.I(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11005__A2 (.I(_03286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10660__A1 (.I(_03286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09323__A2 (.I(_03286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09061__A2 (.I(_03286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07950__I (.I(_03286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08896__A2 (.I(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08768__A2 (.I(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08581__A2 (.I(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08323__A2 (.I(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07951__A2 (.I(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07967__S (.I(_03288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07965__S (.I(_03288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07963__S (.I(_03288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07952__I (.I(_03288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07961__S (.I(_03289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07959__S (.I(_03289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07957__S (.I(_03289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07955__S (.I(_03289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07953__S (.I(_03289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07987__A2 (.I(_03298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07976__I (.I(_03298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07971__I (.I(_03298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07970__I (.I(_03298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07982__A2 (.I(_03299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07980__A2 (.I(_03299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07978__A2 (.I(_03299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07975__A2 (.I(_03299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07973__A2 (.I(_03299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07988__A2 (.I(_03300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07986__A2 (.I(_03300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07984__A2 (.I(_03300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07974__A2 (.I(_03300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07972__A2 (.I(_03300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07985__A2 (.I(_03303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07983__A2 (.I(_03303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07981__A2 (.I(_03303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07979__A2 (.I(_03303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07977__A2 (.I(_03303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10830__A2 (.I(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10387__A2 (.I(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09235__A2 (.I(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08189__A2 (.I(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07990__A2 (.I(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08008__A2 (.I(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07997__I (.I(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07992__I (.I(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07991__I (.I(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08003__A2 (.I(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08001__A2 (.I(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07999__A2 (.I(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07996__A2 (.I(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07994__A2 (.I(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08009__A2 (.I(_03313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08007__A2 (.I(_03313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08005__A2 (.I(_03313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07995__A2 (.I(_03313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07993__A2 (.I(_03313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08006__A2 (.I(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08004__A2 (.I(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08002__A2 (.I(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08000__A2 (.I(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07998__A2 (.I(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08023__A2 (.I(_03324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08021__A2 (.I(_03324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08019__A2 (.I(_03324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08016__A2 (.I(_03324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08014__A2 (.I(_03324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08029__A2 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08027__A2 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08025__A2 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08015__A2 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08013__A2 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08026__A2 (.I(_03328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08024__A2 (.I(_03328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08022__A2 (.I(_03328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08020__A2 (.I(_03328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08018__A2 (.I(_03328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08124__A1 (.I(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08104__A1 (.I(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08083__A1 (.I(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08062__A1 (.I(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08035__A1 (.I(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08048__A2 (.I(_03337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08045__A2 (.I(_03337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08042__A2 (.I(_03337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08038__A2 (.I(_03337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08035__A2 (.I(_03337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08057__A2 (.I(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08054__A2 (.I(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08051__A2 (.I(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08037__A2 (.I(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08034__A2 (.I(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08126__A1 (.I(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08106__A1 (.I(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08085__A1 (.I(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08064__A1 (.I(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08038__A1 (.I(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08129__A1 (.I(_03342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08109__A1 (.I(_03342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08088__A1 (.I(_03342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08067__A1 (.I(_03342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08042__A1 (.I(_03342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08131__A1 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08111__A1 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08090__A1 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08069__A1 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08045__A1 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08133__A1 (.I(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08113__A1 (.I(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08092__A1 (.I(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08071__A1 (.I(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08048__A1 (.I(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08135__A1 (.I(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08115__A1 (.I(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08094__A1 (.I(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08073__A1 (.I(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08051__A1 (.I(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08137__A1 (.I(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08117__A1 (.I(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08096__A1 (.I(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08075__A1 (.I(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08054__A1 (.I(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08139__A1 (.I(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08119__A1 (.I(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08098__A1 (.I(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08077__A1 (.I(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08057__A1 (.I(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08071__A2 (.I(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08069__A2 (.I(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08067__A2 (.I(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08064__A2 (.I(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08062__A2 (.I(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10260__A1 (.I(_03367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10161__A1 (.I(_03367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08896__A1 (.I(_03367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08189__A1 (.I(_03367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08079__A1 (.I(_03367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08092__A2 (.I(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08090__A2 (.I(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08088__A2 (.I(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08085__A2 (.I(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08083__A2 (.I(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08098__A2 (.I(_03370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08096__A2 (.I(_03370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08094__A2 (.I(_03370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08084__A2 (.I(_03370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08082__A2 (.I(_03370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08708__A2 (.I(_03380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08323__A1 (.I(_03380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08269__A1 (.I(_03380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08247__A1 (.I(_03380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08100__A1 (.I(_03380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08119__A2 (.I(_03383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08117__A2 (.I(_03383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08115__A2 (.I(_03383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08105__A2 (.I(_03383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08103__A2 (.I(_03383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08116__A2 (.I(_03386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08114__A2 (.I(_03386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08112__A2 (.I(_03386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08110__A2 (.I(_03386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08108__A2 (.I(_03386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08133__A2 (.I(_03394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08131__A2 (.I(_03394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08129__A2 (.I(_03394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08126__A2 (.I(_03394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08124__A2 (.I(_03394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08139__A2 (.I(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08137__A2 (.I(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08135__A2 (.I(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08125__A2 (.I(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08123__A2 (.I(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08251__A1 (.I(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08231__A1 (.I(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08193__A1 (.I(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08173__A1 (.I(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08145__A1 (.I(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08158__A2 (.I(_03407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08155__A2 (.I(_03407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08152__A2 (.I(_03407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08148__A2 (.I(_03407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08145__A2 (.I(_03407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08167__A2 (.I(_03408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08164__A2 (.I(_03408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08161__A2 (.I(_03408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08147__A2 (.I(_03408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08144__A2 (.I(_03408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08253__A1 (.I(_03410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08233__A1 (.I(_03410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08195__A1 (.I(_03410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08175__A1 (.I(_03410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08148__A1 (.I(_03410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08256__A1 (.I(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08236__A1 (.I(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08198__A1 (.I(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08178__A1 (.I(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08152__A1 (.I(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08258__A1 (.I(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08238__A1 (.I(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08200__A1 (.I(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08180__A1 (.I(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08155__A1 (.I(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08260__A1 (.I(_03417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08240__A1 (.I(_03417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08202__A1 (.I(_03417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08182__A1 (.I(_03417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08158__A1 (.I(_03417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08262__A1 (.I(_03419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08242__A1 (.I(_03419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08204__A1 (.I(_03419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08184__A1 (.I(_03419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08161__A1 (.I(_03419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08264__A1 (.I(_03421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08244__A1 (.I(_03421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08206__A1 (.I(_03421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08186__A1 (.I(_03421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08164__A1 (.I(_03421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08266__A1 (.I(_03423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08246__A1 (.I(_03423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08208__A1 (.I(_03423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08188__A1 (.I(_03423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08167__A1 (.I(_03423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08363__A2 (.I(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08343__A2 (.I(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08303__A2 (.I(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08227__A2 (.I(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08169__A2 (.I(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08188__A2 (.I(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08186__A2 (.I(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08184__A2 (.I(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08174__A2 (.I(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08172__A2 (.I(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08185__A2 (.I(_03431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08183__A2 (.I(_03431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08181__A2 (.I(_03431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08179__A2 (.I(_03431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08177__A2 (.I(_03431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08207__A2 (.I(_03438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08196__I (.I(_03438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08191__I (.I(_03438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08190__I (.I(_03438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08202__A2 (.I(_03439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08200__A2 (.I(_03439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08198__A2 (.I(_03439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08195__A2 (.I(_03439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08193__A2 (.I(_03439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08208__A2 (.I(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08206__A2 (.I(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08204__A2 (.I(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08194__A2 (.I(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08192__A2 (.I(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08225__S (.I(_03450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08223__S (.I(_03450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08221__S (.I(_03450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08210__I (.I(_03450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08219__S (.I(_03451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08217__S (.I(_03451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08215__S (.I(_03451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08213__S (.I(_03451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08211__S (.I(_03451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08245__A2 (.I(_03460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08234__I (.I(_03460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08229__I (.I(_03460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08228__I (.I(_03460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08240__A2 (.I(_03461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08238__A2 (.I(_03461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08236__A2 (.I(_03461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08233__A2 (.I(_03461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08231__A2 (.I(_03461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08246__A2 (.I(_03462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08244__A2 (.I(_03462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08242__A2 (.I(_03462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08232__A2 (.I(_03462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08230__A2 (.I(_03462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08243__A2 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08241__A2 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08239__A2 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08237__A2 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08235__A2 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08265__A2 (.I(_03472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08254__I (.I(_03472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08249__I (.I(_03472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08248__I (.I(_03472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08260__A2 (.I(_03473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08258__A2 (.I(_03473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08256__A2 (.I(_03473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08253__A2 (.I(_03473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08251__A2 (.I(_03473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08266__A2 (.I(_03474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08264__A2 (.I(_03474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08262__A2 (.I(_03474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08252__A2 (.I(_03474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08250__A2 (.I(_03474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08263__A2 (.I(_03477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08261__A2 (.I(_03477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08259__A2 (.I(_03477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08257__A2 (.I(_03477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08255__A2 (.I(_03477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08788__I (.I(_03484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08680__I (.I(_03484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08553__I (.I(_03484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08427__I (.I(_03484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08268__I (.I(_03484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08367__A1 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08347__A1 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08327__A1 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08307__A1 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08273__A1 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08302__A2 (.I(_03488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08298__A2 (.I(_03488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08294__A2 (.I(_03488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08276__A2 (.I(_03488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08272__A2 (.I(_03488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08795__I (.I(_03490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08686__I (.I(_03490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08559__I (.I(_03490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08433__I (.I(_03490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08275__I (.I(_03490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08369__A1 (.I(_03491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08349__A1 (.I(_03491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08329__A1 (.I(_03491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08309__A1 (.I(_03491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08277__A1 (.I(_03491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08798__I (.I(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08689__I (.I(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08562__I (.I(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08436__I (.I(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08279__I (.I(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08372__A1 (.I(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08352__A1 (.I(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08332__A1 (.I(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08312__A1 (.I(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08282__A1 (.I(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08297__A2 (.I(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08293__A2 (.I(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08289__A2 (.I(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08285__A2 (.I(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08281__A2 (.I(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08802__I (.I(_03497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08693__I (.I(_03497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08566__I (.I(_03497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08440__I (.I(_03497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08284__I (.I(_03497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08374__A1 (.I(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08354__A1 (.I(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08334__A1 (.I(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08314__A1 (.I(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08286__A1 (.I(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08805__I (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08696__I (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08569__I (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08443__I (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08288__I (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08376__A1 (.I(_03501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08356__A1 (.I(_03501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08336__A1 (.I(_03501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08316__A1 (.I(_03501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08290__A1 (.I(_03501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08808__I (.I(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08699__I (.I(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08572__I (.I(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08446__I (.I(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08292__I (.I(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08378__A1 (.I(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08358__A1 (.I(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08338__A1 (.I(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08318__A1 (.I(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08294__A1 (.I(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08811__I (.I(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08702__I (.I(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08575__I (.I(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08449__I (.I(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08296__I (.I(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08380__A1 (.I(_03507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08360__A1 (.I(_03507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08340__A1 (.I(_03507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08320__A1 (.I(_03507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08298__A1 (.I(_03507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08814__I (.I(_03509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08705__I (.I(_03509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08578__I (.I(_03509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08452__I (.I(_03509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08300__I (.I(_03509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08382__A1 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08362__A1 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08342__A1 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08322__A1 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08302__A1 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08316__A2 (.I(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08314__A2 (.I(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08312__A2 (.I(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08309__A2 (.I(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08307__A2 (.I(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08322__A2 (.I(_03514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08320__A2 (.I(_03514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08318__A2 (.I(_03514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08308__A2 (.I(_03514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08306__A2 (.I(_03514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08319__A2 (.I(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08317__A2 (.I(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08315__A2 (.I(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08313__A2 (.I(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08311__A2 (.I(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08336__A2 (.I(_03525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08334__A2 (.I(_03525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08332__A2 (.I(_03525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08329__A2 (.I(_03525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08327__A2 (.I(_03525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08342__A2 (.I(_03526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08340__A2 (.I(_03526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08338__A2 (.I(_03526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08328__A2 (.I(_03526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08326__A2 (.I(_03526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08339__A2 (.I(_03529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08337__A2 (.I(_03529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08335__A2 (.I(_03529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08333__A2 (.I(_03529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08331__A2 (.I(_03529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08356__A2 (.I(_03537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08354__A2 (.I(_03537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08352__A2 (.I(_03537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08349__A2 (.I(_03537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08347__A2 (.I(_03537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08362__A2 (.I(_03538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08360__A2 (.I(_03538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08358__A2 (.I(_03538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08348__A2 (.I(_03538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08346__A2 (.I(_03538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08359__A2 (.I(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08357__A2 (.I(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08355__A2 (.I(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08353__A2 (.I(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08351__A2 (.I(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08381__A2 (.I(_03548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08370__I (.I(_03548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08365__I (.I(_03548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08364__I (.I(_03548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08376__A2 (.I(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08374__A2 (.I(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08372__A2 (.I(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08369__A2 (.I(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08367__A2 (.I(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08382__A2 (.I(_03550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08380__A2 (.I(_03550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08378__A2 (.I(_03550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08368__A2 (.I(_03550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08366__A2 (.I(_03550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08379__A2 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08377__A2 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08375__A2 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08373__A2 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08371__A2 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08880__I0 (.I(_03560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08624__I0 (.I(_03560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08497__I0 (.I(_03560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08411__I0 (.I(_03560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08386__I0 (.I(_03560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08407__S (.I(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08404__S (.I(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08401__S (.I(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08385__I (.I(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08882__I0 (.I(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08626__I0 (.I(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08499__I0 (.I(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08413__I0 (.I(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08389__I0 (.I(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08884__I0 (.I(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08628__I0 (.I(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08501__I0 (.I(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08415__I0 (.I(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08392__I0 (.I(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08886__I0 (.I(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08630__I0 (.I(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08503__I0 (.I(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08417__I0 (.I(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08395__I0 (.I(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08888__I0 (.I(_03570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08632__I0 (.I(_03570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08505__I0 (.I(_03570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08419__I0 (.I(_03570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08398__I0 (.I(_03570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08890__I0 (.I(_03572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08634__I0 (.I(_03572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08507__I0 (.I(_03572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08421__I0 (.I(_03572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08401__I0 (.I(_03572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08892__I0 (.I(_03574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08636__I0 (.I(_03574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08509__I0 (.I(_03574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08423__I0 (.I(_03574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08404__I0 (.I(_03574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08894__I0 (.I(_03576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08638__I0 (.I(_03576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08511__I0 (.I(_03576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08425__I0 (.I(_03576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08407__I0 (.I(_03576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08425__S (.I(_03578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08423__S (.I(_03578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08421__S (.I(_03578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08410__I (.I(_03578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08419__S (.I(_03579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08417__S (.I(_03579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08415__S (.I(_03579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08413__S (.I(_03579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08411__S (.I(_03579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08537__A1 (.I(_03588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08517__A1 (.I(_03588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08479__A1 (.I(_03588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08459__A1 (.I(_03588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08432__A1 (.I(_03588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08453__A2 (.I(_03589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08437__I (.I(_03589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08430__I (.I(_03589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08429__I (.I(_03589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08445__A2 (.I(_03590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08442__A2 (.I(_03590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08439__A2 (.I(_03590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08435__A2 (.I(_03590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08432__A2 (.I(_03590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08454__A2 (.I(_03591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08451__A2 (.I(_03591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08448__A2 (.I(_03591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08434__A2 (.I(_03591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08431__A2 (.I(_03591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08539__A1 (.I(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08519__A1 (.I(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08481__A1 (.I(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08461__A1 (.I(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08435__A1 (.I(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08542__A1 (.I(_03595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08522__A1 (.I(_03595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08484__A1 (.I(_03595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08464__A1 (.I(_03595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08439__A1 (.I(_03595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08450__A2 (.I(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08447__A2 (.I(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08444__A2 (.I(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08441__A2 (.I(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08438__A2 (.I(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08544__A1 (.I(_03598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08524__A1 (.I(_03598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08486__A1 (.I(_03598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08466__A1 (.I(_03598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08442__A1 (.I(_03598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08546__A1 (.I(_03600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08526__A1 (.I(_03600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08488__A1 (.I(_03600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08468__A1 (.I(_03600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08445__A1 (.I(_03600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08548__A1 (.I(_03602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08528__A1 (.I(_03602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08490__A1 (.I(_03602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08470__A1 (.I(_03602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08448__A1 (.I(_03602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08550__A1 (.I(_03604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08530__A1 (.I(_03604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08492__A1 (.I(_03604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08472__A1 (.I(_03604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08451__A1 (.I(_03604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08552__A1 (.I(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08532__A1 (.I(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08494__A1 (.I(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08474__A1 (.I(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08454__A1 (.I(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08473__A2 (.I(_03608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08462__I (.I(_03608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08457__I (.I(_03608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08456__I (.I(_03608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08468__A2 (.I(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08466__A2 (.I(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08464__A2 (.I(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08461__A2 (.I(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08459__A2 (.I(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08474__A2 (.I(_03610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08472__A2 (.I(_03610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08470__A2 (.I(_03610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08460__A2 (.I(_03610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08458__A2 (.I(_03610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08471__A2 (.I(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08469__A2 (.I(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08467__A2 (.I(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08465__A2 (.I(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08463__A2 (.I(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08493__A2 (.I(_03620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08482__I (.I(_03620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08477__I (.I(_03620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08476__I (.I(_03620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08488__A2 (.I(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08486__A2 (.I(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08484__A2 (.I(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08481__A2 (.I(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08479__A2 (.I(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08494__A2 (.I(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08492__A2 (.I(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08490__A2 (.I(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08480__A2 (.I(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08478__A2 (.I(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08491__A2 (.I(_03625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08489__A2 (.I(_03625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08487__A2 (.I(_03625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08485__A2 (.I(_03625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08483__A2 (.I(_03625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08511__S (.I(_03632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08509__S (.I(_03632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08507__S (.I(_03632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08496__I (.I(_03632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08505__S (.I(_03633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08503__S (.I(_03633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08501__S (.I(_03633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08499__S (.I(_03633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08497__S (.I(_03633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08526__A2 (.I(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08524__A2 (.I(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08522__A2 (.I(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08519__A2 (.I(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08517__A2 (.I(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08532__A2 (.I(_03644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08530__A2 (.I(_03644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08528__A2 (.I(_03644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08518__A2 (.I(_03644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08516__A2 (.I(_03644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08529__A2 (.I(_03647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08527__A2 (.I(_03647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08525__A2 (.I(_03647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08523__A2 (.I(_03647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08521__A2 (.I(_03647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08546__A2 (.I(_03655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08544__A2 (.I(_03655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08542__A2 (.I(_03655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08539__A2 (.I(_03655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08537__A2 (.I(_03655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08552__A2 (.I(_03656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08550__A2 (.I(_03656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08548__A2 (.I(_03656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08538__A2 (.I(_03656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08536__A2 (.I(_03656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08549__A2 (.I(_03659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08547__A2 (.I(_03659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08545__A2 (.I(_03659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08543__A2 (.I(_03659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08541__A2 (.I(_03659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08664__A1 (.I(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08644__A1 (.I(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08606__A1 (.I(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08585__A1 (.I(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08558__A1 (.I(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08666__A1 (.I(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08646__A1 (.I(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08608__A1 (.I(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08587__A1 (.I(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08561__A1 (.I(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08669__A1 (.I(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08649__A1 (.I(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08611__A1 (.I(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08590__A1 (.I(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08565__A1 (.I(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08576__A2 (.I(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08573__A2 (.I(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08570__A2 (.I(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08567__A2 (.I(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08564__A2 (.I(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08671__A1 (.I(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08651__A1 (.I(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08613__A1 (.I(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08592__A1 (.I(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08568__A1 (.I(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08673__A1 (.I(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08653__A1 (.I(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08615__A1 (.I(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08594__A1 (.I(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08571__A1 (.I(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08675__A1 (.I(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08655__A1 (.I(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08617__A1 (.I(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08596__A1 (.I(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08574__A1 (.I(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08677__A1 (.I(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08657__A1 (.I(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08619__A1 (.I(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08598__A1 (.I(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08577__A1 (.I(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08679__A1 (.I(_03684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08659__A1 (.I(_03684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08621__A1 (.I(_03684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08600__A1 (.I(_03684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08580__A1 (.I(_03684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08600__A2 (.I(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08598__A2 (.I(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08596__A2 (.I(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08586__A2 (.I(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08584__A2 (.I(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08597__A2 (.I(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08595__A2 (.I(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08593__A2 (.I(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08591__A2 (.I(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08589__A2 (.I(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08748__A2 (.I(_03698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08728__A2 (.I(_03698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08681__A2 (.I(_03698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08640__A2 (.I(_03698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08602__A2 (.I(_03698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08615__A2 (.I(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08613__A2 (.I(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08611__A2 (.I(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08608__A2 (.I(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08606__A2 (.I(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08621__A2 (.I(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08619__A2 (.I(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08617__A2 (.I(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08607__A2 (.I(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08605__A2 (.I(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08618__A2 (.I(_03704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08616__A2 (.I(_03704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08614__A2 (.I(_03704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08612__A2 (.I(_03704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08610__A2 (.I(_03704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08638__S (.I(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08636__S (.I(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08634__S (.I(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08623__I (.I(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08632__S (.I(_03712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08630__S (.I(_03712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08628__S (.I(_03712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08626__S (.I(_03712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08624__S (.I(_03712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08656__A2 (.I(_03726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08654__A2 (.I(_03726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08652__A2 (.I(_03726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08650__A2 (.I(_03726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08648__A2 (.I(_03726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08673__A2 (.I(_03734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08671__A2 (.I(_03734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08669__A2 (.I(_03734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08666__A2 (.I(_03734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08664__A2 (.I(_03734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08772__A1 (.I(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08752__A1 (.I(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08732__A1 (.I(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08712__A1 (.I(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08685__A1 (.I(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08698__A2 (.I(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08695__A2 (.I(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08692__A2 (.I(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08688__A2 (.I(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08685__A2 (.I(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08707__A2 (.I(_03748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08704__A2 (.I(_03748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08701__A2 (.I(_03748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08687__A2 (.I(_03748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08684__A2 (.I(_03748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08774__A1 (.I(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08754__A1 (.I(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08734__A1 (.I(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08714__A1 (.I(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08688__A1 (.I(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08777__A1 (.I(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08757__A1 (.I(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08737__A1 (.I(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08717__A1 (.I(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08692__A1 (.I(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08703__A2 (.I(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08700__A2 (.I(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08697__A2 (.I(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08694__A2 (.I(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08691__A2 (.I(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08779__A1 (.I(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08759__A1 (.I(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08739__A1 (.I(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08719__A1 (.I(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08695__A1 (.I(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08781__A1 (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08761__A1 (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08741__A1 (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08721__A1 (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08698__A1 (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08783__A1 (.I(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08763__A1 (.I(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08743__A1 (.I(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08723__A1 (.I(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08701__A1 (.I(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08785__A1 (.I(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08765__A1 (.I(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08745__A1 (.I(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08725__A1 (.I(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08704__A1 (.I(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08787__A1 (.I(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08767__A1 (.I(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08747__A1 (.I(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08727__A1 (.I(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08707__A1 (.I(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08727__A2 (.I(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08725__A2 (.I(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08723__A2 (.I(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08713__A2 (.I(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08711__A2 (.I(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08746__A2 (.I(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08735__I (.I(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08730__I (.I(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08729__I (.I(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08741__A2 (.I(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08739__A2 (.I(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08737__A2 (.I(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08734__A2 (.I(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08732__A2 (.I(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08744__A2 (.I(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08742__A2 (.I(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08740__A2 (.I(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08738__A2 (.I(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08736__A2 (.I(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08766__A2 (.I(_03789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08755__I (.I(_03789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08750__I (.I(_03789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08749__I (.I(_03789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08761__A2 (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08759__A2 (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08757__A2 (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08754__A2 (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08752__A2 (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08767__A2 (.I(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08765__A2 (.I(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08763__A2 (.I(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08753__A2 (.I(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08751__A2 (.I(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08764__A2 (.I(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08762__A2 (.I(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08760__A2 (.I(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08758__A2 (.I(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08756__A2 (.I(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08786__A2 (.I(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08775__I (.I(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08770__I (.I(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08769__I (.I(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08781__A2 (.I(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08779__A2 (.I(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08777__A2 (.I(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08774__A2 (.I(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08772__A2 (.I(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08787__A2 (.I(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08785__A2 (.I(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08783__A2 (.I(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08773__A2 (.I(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08771__A2 (.I(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08784__A2 (.I(_03806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08782__A2 (.I(_03806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08780__A2 (.I(_03806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08778__A2 (.I(_03806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08776__A2 (.I(_03806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08900__A1 (.I(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08861__A1 (.I(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08841__A1 (.I(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08821__A1 (.I(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08794__A1 (.I(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08918__A2 (.I(_03814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08857__A2 (.I(_03814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08837__A2 (.I(_03814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08817__A2 (.I(_03814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08790__A2 (.I(_03814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08815__A2 (.I(_03815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08799__I (.I(_03815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08792__I (.I(_03815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08791__I (.I(_03815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08807__A2 (.I(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08804__A2 (.I(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08801__A2 (.I(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08797__A2 (.I(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08794__A2 (.I(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08816__A2 (.I(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08813__A2 (.I(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08810__A2 (.I(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08796__A2 (.I(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08793__A2 (.I(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08902__A1 (.I(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08863__A1 (.I(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08843__A1 (.I(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08823__A1 (.I(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08797__A1 (.I(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08905__A1 (.I(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08866__A1 (.I(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08846__A1 (.I(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08826__A1 (.I(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08801__A1 (.I(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08812__A2 (.I(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08809__A2 (.I(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08806__A2 (.I(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08803__A2 (.I(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08800__A2 (.I(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08907__A1 (.I(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08868__A1 (.I(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08848__A1 (.I(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08828__A1 (.I(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08804__A1 (.I(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08909__A1 (.I(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08870__A1 (.I(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08850__A1 (.I(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08830__A1 (.I(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08807__A1 (.I(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08911__A1 (.I(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08872__A1 (.I(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08852__A1 (.I(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08832__A1 (.I(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08810__A1 (.I(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08913__A1 (.I(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08874__A1 (.I(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08854__A1 (.I(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08834__A1 (.I(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08813__A1 (.I(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08915__A1 (.I(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08876__A1 (.I(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08856__A1 (.I(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08836__A1 (.I(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08816__A1 (.I(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08835__A2 (.I(_03834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08824__I (.I(_03834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08819__I (.I(_03834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08818__I (.I(_03834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08830__A2 (.I(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08828__A2 (.I(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08826__A2 (.I(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08823__A2 (.I(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08821__A2 (.I(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08836__A2 (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08834__A2 (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08832__A2 (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08822__A2 (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08820__A2 (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08833__A2 (.I(_03839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08831__A2 (.I(_03839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08829__A2 (.I(_03839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08827__A2 (.I(_03839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08825__A2 (.I(_03839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08855__A2 (.I(_03846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08844__I (.I(_03846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08839__I (.I(_03846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08838__I (.I(_03846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08850__A2 (.I(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08848__A2 (.I(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08846__A2 (.I(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08843__A2 (.I(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08841__A2 (.I(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08856__A2 (.I(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08854__A2 (.I(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08852__A2 (.I(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08842__A2 (.I(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08840__A2 (.I(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08853__A2 (.I(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08851__A2 (.I(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08849__A2 (.I(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08847__A2 (.I(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08845__A2 (.I(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08875__A2 (.I(_03858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08864__I (.I(_03858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08859__I (.I(_03858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08858__I (.I(_03858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08870__A2 (.I(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08868__A2 (.I(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08866__A2 (.I(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08863__A2 (.I(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08861__A2 (.I(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08876__A2 (.I(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08874__A2 (.I(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08872__A2 (.I(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08862__A2 (.I(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08860__A2 (.I(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08873__A2 (.I(_03863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08871__A2 (.I(_03863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08869__A2 (.I(_03863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08867__A2 (.I(_03863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08865__A2 (.I(_03863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08894__S (.I(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08892__S (.I(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08890__S (.I(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08879__I (.I(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08888__S (.I(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08886__S (.I(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08884__S (.I(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08882__S (.I(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08880__S (.I(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08914__A2 (.I(_03881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08903__I (.I(_03881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08898__I (.I(_03881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08897__I (.I(_03881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08909__A2 (.I(_03882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08907__A2 (.I(_03882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08905__A2 (.I(_03882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08902__A2 (.I(_03882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08900__A2 (.I(_03882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08915__A2 (.I(_03883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08913__A2 (.I(_03883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08911__A2 (.I(_03883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08901__A2 (.I(_03883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08899__A2 (.I(_03883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08912__A2 (.I(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08910__A2 (.I(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08908__A2 (.I(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08906__A2 (.I(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08904__A2 (.I(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09448__I (.I(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09295__I (.I(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09167__I (.I(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09032__I (.I(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08917__I (.I(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09016__A1 (.I(_03894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08996__A1 (.I(_03894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08976__A1 (.I(_03894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08956__A1 (.I(_03894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08922__A1 (.I(_03894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08950__A2 (.I(_03895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08929__I (.I(_03895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08920__I (.I(_03895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08919__I (.I(_03895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08939__A2 (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08935__A2 (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08931__A2 (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08926__A2 (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08922__A2 (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08951__A2 (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08947__A2 (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08943__A2 (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08925__A2 (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08921__A2 (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09454__I (.I(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09301__I (.I(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09173__I (.I(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09039__I (.I(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08924__I (.I(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09018__A1 (.I(_03900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08998__A1 (.I(_03900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08978__A1 (.I(_03900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08958__A1 (.I(_03900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08926__A1 (.I(_03900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09457__I (.I(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09304__I (.I(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09176__I (.I(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09042__I (.I(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08928__I (.I(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09021__A1 (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09001__A1 (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08981__A1 (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08961__A1 (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08931__A1 (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08946__A2 (.I(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08942__A2 (.I(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08938__A2 (.I(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08934__A2 (.I(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08930__A2 (.I(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09461__I (.I(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09308__I (.I(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09180__I (.I(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09046__I (.I(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08933__I (.I(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09023__A1 (.I(_03907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09003__A1 (.I(_03907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08983__A1 (.I(_03907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08963__A1 (.I(_03907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08935__A1 (.I(_03907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09464__I (.I(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09311__I (.I(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09183__I (.I(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09049__I (.I(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08937__I (.I(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09025__A1 (.I(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09005__A1 (.I(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08985__A1 (.I(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08965__A1 (.I(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08939__A1 (.I(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09467__I (.I(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09314__I (.I(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09186__I (.I(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09052__I (.I(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08941__I (.I(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09027__A1 (.I(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09007__A1 (.I(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08987__A1 (.I(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08967__A1 (.I(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08943__A1 (.I(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09470__I (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09317__I (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09189__I (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09055__I (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08945__I (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09029__A1 (.I(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09009__A1 (.I(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08989__A1 (.I(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08969__A1 (.I(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08947__A1 (.I(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09473__I (.I(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09320__I (.I(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09192__I (.I(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09058__I (.I(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08949__I (.I(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09031__A1 (.I(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09011__A1 (.I(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08991__A1 (.I(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08971__A1 (.I(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08951__A1 (.I(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08970__A2 (.I(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08959__I (.I(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08954__I (.I(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08953__I (.I(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08965__A2 (.I(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08963__A2 (.I(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08961__A2 (.I(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08958__A2 (.I(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08956__A2 (.I(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08971__A2 (.I(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08969__A2 (.I(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08967__A2 (.I(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08957__A2 (.I(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08955__A2 (.I(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08968__A2 (.I(_03926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08966__A2 (.I(_03926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08964__A2 (.I(_03926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08962__A2 (.I(_03926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08960__A2 (.I(_03926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08990__A2 (.I(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08979__I (.I(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08974__I (.I(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08973__I (.I(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08985__A2 (.I(_03934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08983__A2 (.I(_03934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08981__A2 (.I(_03934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08978__A2 (.I(_03934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08976__A2 (.I(_03934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08991__A2 (.I(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08989__A2 (.I(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08987__A2 (.I(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08977__A2 (.I(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08975__A2 (.I(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08988__A2 (.I(_03938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08986__A2 (.I(_03938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08984__A2 (.I(_03938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08982__A2 (.I(_03938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08980__A2 (.I(_03938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09010__A2 (.I(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08999__I (.I(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08994__I (.I(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08993__I (.I(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09005__A2 (.I(_03946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09003__A2 (.I(_03946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09001__A2 (.I(_03946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08998__A2 (.I(_03946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08996__A2 (.I(_03946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09011__A2 (.I(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09009__A2 (.I(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09007__A2 (.I(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08997__A2 (.I(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08995__A2 (.I(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09008__A2 (.I(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09006__A2 (.I(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09004__A2 (.I(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09002__A2 (.I(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09000__A2 (.I(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09030__A2 (.I(_03957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09019__I (.I(_03957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09014__I (.I(_03957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09013__I (.I(_03957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09025__A2 (.I(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09023__A2 (.I(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09021__A2 (.I(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09018__A2 (.I(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09016__A2 (.I(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09031__A2 (.I(_03959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09029__A2 (.I(_03959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09027__A2 (.I(_03959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09017__A2 (.I(_03959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09015__A2 (.I(_03959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09028__A2 (.I(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09026__A2 (.I(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09024__A2 (.I(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09022__A2 (.I(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09020__A2 (.I(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09151__A1 (.I(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09105__A1 (.I(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09085__A1 (.I(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09065__A1 (.I(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09038__A1 (.I(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09407__A2 (.I(_03970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09343__A2 (.I(_03970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09296__A2 (.I(_03970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09275__A2 (.I(_03970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09034__A2 (.I(_03970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09060__A2 (.I(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09057__A2 (.I(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09054__A2 (.I(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09040__A2 (.I(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09037__A2 (.I(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09153__A1 (.I(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09107__A1 (.I(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09087__A1 (.I(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09067__A1 (.I(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09041__A1 (.I(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09156__A1 (.I(_03977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09110__A1 (.I(_03977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09090__A1 (.I(_03977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09070__A1 (.I(_03977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09045__A1 (.I(_03977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09056__A2 (.I(_03978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09053__A2 (.I(_03978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09050__A2 (.I(_03978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09047__A2 (.I(_03978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09044__A2 (.I(_03978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09158__A1 (.I(_03980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09112__A1 (.I(_03980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09092__A1 (.I(_03980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09072__A1 (.I(_03980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09048__A1 (.I(_03980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09160__A1 (.I(_03982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09114__A1 (.I(_03982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09094__A1 (.I(_03982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09074__A1 (.I(_03982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09051__A1 (.I(_03982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09162__A1 (.I(_03984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09116__A1 (.I(_03984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09096__A1 (.I(_03984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09076__A1 (.I(_03984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09054__A1 (.I(_03984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09164__A1 (.I(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09118__A1 (.I(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09098__A1 (.I(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09078__A1 (.I(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09057__A1 (.I(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09166__A1 (.I(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09120__A1 (.I(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09100__A1 (.I(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09080__A1 (.I(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09060__A1 (.I(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09079__A2 (.I(_03990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09068__I (.I(_03990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09063__I (.I(_03990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09062__I (.I(_03990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09077__A2 (.I(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09075__A2 (.I(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09073__A2 (.I(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09071__A2 (.I(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09069__A2 (.I(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09100__A2 (.I(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09098__A2 (.I(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09096__A2 (.I(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09086__A2 (.I(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09084__A2 (.I(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09097__A2 (.I(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09095__A2 (.I(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09093__A2 (.I(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09091__A2 (.I(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09089__A2 (.I(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09117__A2 (.I(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09115__A2 (.I(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09113__A2 (.I(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09111__A2 (.I(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09109__A2 (.I(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11105__A1 (.I(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11085__A1 (.I(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10122__A1 (.I(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09136__A2 (.I(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09122__A1 (.I(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11111__A3 (.I(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09516__B (.I(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09133__A1 (.I(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09131__A1 (.I(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09130__A1 (.I(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11317__A1 (.I(_04032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11113__B (.I(_04032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09142__A1 (.I(_04032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09140__C (.I(_04032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09130__B (.I(_04032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11111__A2 (.I(_04034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09517__A2 (.I(_04034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09516__A2 (.I(_04034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09210__A1 (.I(_04034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09134__A1 (.I(_04034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09165__A2 (.I(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09154__I (.I(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09149__I (.I(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09148__I (.I(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09163__A2 (.I(_04049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09161__A2 (.I(_04049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09159__A2 (.I(_04049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09157__A2 (.I(_04049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09155__A2 (.I(_04049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09279__A1 (.I(_04056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09259__A1 (.I(_04056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09239__A1 (.I(_04056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09219__A1 (.I(_04056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09172__A1 (.I(_04056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09193__A2 (.I(_04057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09177__I (.I(_04057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09170__I (.I(_04057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09169__I (.I(_04057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09185__A2 (.I(_04058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09182__A2 (.I(_04058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09179__A2 (.I(_04058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09175__A2 (.I(_04058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09172__A2 (.I(_04058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09194__A2 (.I(_04059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09191__A2 (.I(_04059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09188__A2 (.I(_04059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09174__A2 (.I(_04059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09171__A2 (.I(_04059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09281__A1 (.I(_04061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09261__A1 (.I(_04061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09241__A1 (.I(_04061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09221__A1 (.I(_04061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09175__A1 (.I(_04061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09284__A1 (.I(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09264__A1 (.I(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09244__A1 (.I(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09224__A1 (.I(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09179__A1 (.I(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09190__A2 (.I(_04064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09187__A2 (.I(_04064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09184__A2 (.I(_04064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09181__A2 (.I(_04064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09178__A2 (.I(_04064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09286__A1 (.I(_04066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09266__A1 (.I(_04066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09246__A1 (.I(_04066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09226__A1 (.I(_04066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09182__A1 (.I(_04066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09288__A1 (.I(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09268__A1 (.I(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09248__A1 (.I(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09228__A1 (.I(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09185__A1 (.I(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09290__A1 (.I(_04070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09270__A1 (.I(_04070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09250__A1 (.I(_04070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09230__A1 (.I(_04070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09188__A1 (.I(_04070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09292__A1 (.I(_04072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09272__A1 (.I(_04072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09252__A1 (.I(_04072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09232__A1 (.I(_04072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09191__A1 (.I(_04072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09294__A1 (.I(_04074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09274__A1 (.I(_04074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09254__A1 (.I(_04074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09234__A1 (.I(_04074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09194__A1 (.I(_04074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10830__A1 (.I(_04091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10531__A1 (.I(_04091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10511__A1 (.I(_04091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10423__A1 (.I(_04091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09215__A1 (.I(_04091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09233__A2 (.I(_04092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09222__I (.I(_04092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09217__I (.I(_04092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09216__I (.I(_04092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09231__A2 (.I(_04097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09229__A2 (.I(_04097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09227__A2 (.I(_04097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09225__A2 (.I(_04097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09223__A2 (.I(_04097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09253__A2 (.I(_04104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09242__I (.I(_04104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09237__I (.I(_04104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09236__I (.I(_04104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09248__A2 (.I(_04105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09246__A2 (.I(_04105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09244__A2 (.I(_04105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09241__A2 (.I(_04105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09239__A2 (.I(_04105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09254__A2 (.I(_04106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09252__A2 (.I(_04106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09250__A2 (.I(_04106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09240__A2 (.I(_04106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09238__A2 (.I(_04106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09251__A2 (.I(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09249__A2 (.I(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09247__A2 (.I(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09245__A2 (.I(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09243__A2 (.I(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09288__A2 (.I(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09286__A2 (.I(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09284__A2 (.I(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09281__A2 (.I(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09279__A2 (.I(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09432__A1 (.I(_04140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09411__A1 (.I(_04140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09347__A1 (.I(_04140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09327__A1 (.I(_04140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09300__A1 (.I(_04140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09321__A2 (.I(_04141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09305__I (.I(_04141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09298__I (.I(_04141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09297__I (.I(_04141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09313__A2 (.I(_04142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09310__A2 (.I(_04142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09307__A2 (.I(_04142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09303__A2 (.I(_04142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09300__A2 (.I(_04142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09322__A2 (.I(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09319__A2 (.I(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09316__A2 (.I(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09302__A2 (.I(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09299__A2 (.I(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09434__A1 (.I(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09413__A1 (.I(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09349__A1 (.I(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09329__A1 (.I(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09303__A1 (.I(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09437__A1 (.I(_04147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09416__A1 (.I(_04147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09352__A1 (.I(_04147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09332__A1 (.I(_04147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09307__A1 (.I(_04147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09439__A1 (.I(_04150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09418__A1 (.I(_04150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09354__A1 (.I(_04150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09334__A1 (.I(_04150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09310__A1 (.I(_04150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09441__A1 (.I(_04152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09420__A1 (.I(_04152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09356__A1 (.I(_04152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09336__A1 (.I(_04152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09313__A1 (.I(_04152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09443__A1 (.I(_04154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09422__A1 (.I(_04154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09358__A1 (.I(_04154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09338__A1 (.I(_04154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09316__A1 (.I(_04154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09445__A1 (.I(_04156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09424__A1 (.I(_04156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09360__A1 (.I(_04156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09340__A1 (.I(_04156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09319__A1 (.I(_04156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09447__A1 (.I(_04158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09426__A1 (.I(_04158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09362__A1 (.I(_04158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09342__A1 (.I(_04158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09322__A1 (.I(_04158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09341__A2 (.I(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09330__I (.I(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09325__I (.I(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09324__I (.I(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09336__A2 (.I(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09334__A2 (.I(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09332__A2 (.I(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09329__A2 (.I(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09327__A2 (.I(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09339__A2 (.I(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09337__A2 (.I(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09335__A2 (.I(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09333__A2 (.I(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09331__A2 (.I(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09356__A2 (.I(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09354__A2 (.I(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09352__A2 (.I(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09349__A2 (.I(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09347__A2 (.I(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09362__A2 (.I(_04174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09360__A2 (.I(_04174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09358__A2 (.I(_04174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09348__A2 (.I(_04174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09346__A2 (.I(_04174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09359__A2 (.I(_04177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09357__A2 (.I(_04177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09355__A2 (.I(_04177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09353__A2 (.I(_04177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09351__A2 (.I(_04177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10941__I0 (.I(_04184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10407__I0 (.I(_04184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10389__I0 (.I(_04184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09391__I0 (.I(_04184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09366__I0 (.I(_04184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09387__S (.I(_04185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09384__S (.I(_04185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09381__S (.I(_04185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09365__I (.I(_04185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09378__S (.I(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09375__S (.I(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09372__S (.I(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09369__S (.I(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09366__S (.I(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10943__I0 (.I(_04188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10409__I0 (.I(_04188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10391__I0 (.I(_04188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09393__I0 (.I(_04188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09369__I0 (.I(_04188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10945__I0 (.I(_04190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10411__I0 (.I(_04190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10393__I0 (.I(_04190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09395__I0 (.I(_04190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09372__I0 (.I(_04190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10947__I0 (.I(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10413__I0 (.I(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10395__I0 (.I(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09397__I0 (.I(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09375__I0 (.I(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10949__I0 (.I(_04194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10415__I0 (.I(_04194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10397__I0 (.I(_04194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09399__I0 (.I(_04194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09378__I0 (.I(_04194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09405__S (.I(_04202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09403__S (.I(_04202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09401__S (.I(_04202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09390__I (.I(_04202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09399__S (.I(_04203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09397__S (.I(_04203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09395__S (.I(_04203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09393__S (.I(_04203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09391__S (.I(_04203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09873__A2 (.I(_04224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09650__A2 (.I(_04224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09476__A2 (.I(_04224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09449__A2 (.I(_04224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09428__A2 (.I(_04224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09446__A2 (.I(_04225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09435__I (.I(_04225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09430__I (.I(_04225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09429__I (.I(_04225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09441__A2 (.I(_04226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09439__A2 (.I(_04226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09437__A2 (.I(_04226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09434__A2 (.I(_04226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09432__A2 (.I(_04226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09447__A2 (.I(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09445__A2 (.I(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09443__A2 (.I(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09433__A2 (.I(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09431__A2 (.I(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09444__A2 (.I(_04230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09442__A2 (.I(_04230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09440__A2 (.I(_04230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09438__A2 (.I(_04230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09436__A2 (.I(_04230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09877__A1 (.I(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09654__A1 (.I(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09500__A1 (.I(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09480__A1 (.I(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09453__A1 (.I(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09466__A2 (.I(_04239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09463__A2 (.I(_04239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09460__A2 (.I(_04239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09456__A2 (.I(_04239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09453__A2 (.I(_04239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09475__A2 (.I(_04240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09472__A2 (.I(_04240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09469__A2 (.I(_04240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09455__A2 (.I(_04240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09452__A2 (.I(_04240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09879__A1 (.I(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09656__A1 (.I(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09502__A1 (.I(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09482__A1 (.I(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09456__A1 (.I(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09882__A1 (.I(_04244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09659__A1 (.I(_04244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09505__A1 (.I(_04244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09485__A1 (.I(_04244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09460__A1 (.I(_04244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09471__A2 (.I(_04245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09468__A2 (.I(_04245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09465__A2 (.I(_04245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09462__A2 (.I(_04245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09459__A2 (.I(_04245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09884__A1 (.I(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09661__A1 (.I(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09507__A1 (.I(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09487__A1 (.I(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09463__A1 (.I(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09886__A1 (.I(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09663__A1 (.I(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09509__A1 (.I(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09489__A1 (.I(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09466__A1 (.I(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09888__A1 (.I(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09665__A1 (.I(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09511__A1 (.I(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09491__A1 (.I(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09469__A1 (.I(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09890__A1 (.I(_04253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09667__A1 (.I(_04253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09513__A1 (.I(_04253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09493__A1 (.I(_04253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09472__A1 (.I(_04253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09892__A1 (.I(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09669__A1 (.I(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09515__A1 (.I(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09495__A1 (.I(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09475__A1 (.I(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09489__A2 (.I(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09487__A2 (.I(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09485__A2 (.I(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09482__A2 (.I(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09480__A2 (.I(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09492__A2 (.I(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09490__A2 (.I(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09488__A2 (.I(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09486__A2 (.I(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09484__A2 (.I(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09515__A2 (.I(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09513__A2 (.I(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09511__A2 (.I(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09501__A2 (.I(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09499__A2 (.I(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09557__A2 (.I(_04284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09529__A2 (.I(_04284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09520__I (.I(_04284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09631__A2 (.I(_04285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09552__B (.I(_04285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09543__A1 (.I(_04285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09535__A1 (.I(_04285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09523__A1 (.I(_04285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09637__A2 (.I(_04293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09625__A2 (.I(_04293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09622__A2 (.I(_04293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09617__A2 (.I(_04293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09531__A2 (.I(_04293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09613__I (.I(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09591__I (.I(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09573__I (.I(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09560__I (.I(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09530__I (.I(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09640__B1 (.I(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09632__B1 (.I(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09628__A2 (.I(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09565__A2 (.I(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09531__B1 (.I(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10108__A2 (.I(_04310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09700__A2 (.I(_04310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09554__A1 (.I(_04310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09619__A2 (.I(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09595__I (.I(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09577__I (.I(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09553__B (.I(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09550__I (.I(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09627__A2 (.I(_04312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09574__A2 (.I(_04312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09564__A2 (.I(_04312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09562__A2 (.I(_04312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09554__A2 (.I(_04312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09603__I (.I(_04318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09583__I (.I(_04318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09568__I (.I(_04318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09558__I (.I(_04318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09636__A2 (.I(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09628__B1 (.I(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09624__A2 (.I(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09565__B1 (.I(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09559__C (.I(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09619__B1 (.I(_04321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09607__B1 (.I(_04321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09598__B1 (.I(_04321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09569__B1 (.I(_04321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09561__I (.I(_04321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09649__A2 (.I(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09647__A2 (.I(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09644__A2 (.I(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09635__A2 (.I(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09562__B1 (.I(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09640__A2 (.I(_04326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09632__A2 (.I(_04326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09607__A2 (.I(_04326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09598__A2 (.I(_04326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09569__A2 (.I(_04326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09619__C1 (.I(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09607__C1 (.I(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09598__C1 (.I(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09571__I (.I(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09569__C1 (.I(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09647__B1 (.I(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09644__B1 (.I(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09580__A2 (.I(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09576__A2 (.I(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09572__A2 (.I(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09588__B1 (.I(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09585__B1 (.I(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09581__B1 (.I(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09578__B1 (.I(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09574__B1 (.I(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09592__A2 (.I(_04334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09588__A2 (.I(_04334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09585__A2 (.I(_04334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09581__A2 (.I(_04334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09578__A2 (.I(_04334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09600__A2 (.I(_04338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09594__A2 (.I(_04338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09590__A2 (.I(_04338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09587__A2 (.I(_04338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09584__A2 (.I(_04338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09610__B1 (.I(_04344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09605__B1 (.I(_04344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09601__B1 (.I(_04344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09596__B1 (.I(_04344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09592__B1 (.I(_04344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09614__A2 (.I(_04347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09610__A2 (.I(_04347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09605__A2 (.I(_04347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09601__A2 (.I(_04347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09596__A2 (.I(_04347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09621__A2 (.I(_04352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09616__A2 (.I(_04352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09612__A2 (.I(_04352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09609__A2 (.I(_04352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09604__A2 (.I(_04352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09637__B1 (.I(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09625__B1 (.I(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09622__B1 (.I(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09617__B1 (.I(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09614__B1 (.I(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09663__A2 (.I(_04384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09661__A2 (.I(_04384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09659__A2 (.I(_04384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09656__A2 (.I(_04384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09654__A2 (.I(_04384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09669__A2 (.I(_04385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09667__A2 (.I(_04385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09665__A2 (.I(_04385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09655__A2 (.I(_04385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09653__A2 (.I(_04385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09666__A2 (.I(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09664__A2 (.I(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09662__A2 (.I(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09660__A2 (.I(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09658__A2 (.I(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10103__A2 (.I(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10018__B2 (.I(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09818__C (.I(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09794__A2 (.I(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09671__I (.I(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09841__A2 (.I(_04396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09825__A2 (.I(_04396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09819__A2 (.I(_04396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09812__A2 (.I(_04396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09738__A2 (.I(_04396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10110__A1 (.I(_04397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09975__A1 (.I(_04397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09929__A1 (.I(_04397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09856__I (.I(_04397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09673__I (.I(_04397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10454__A1 (.I(_04398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09921__A2 (.I(_04398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09872__A2 (.I(_04398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09858__A2 (.I(_04398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09737__A1 (.I(_04398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09908__A1 (.I(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09782__I (.I(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09678__A1 (.I(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09909__A1 (.I(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09783__I (.I(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09678__A2 (.I(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10460__A1 (.I(_04401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10088__A1 (.I(_04401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09992__A1 (.I(_04401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09678__A3 (.I(_04401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10033__A1 (.I(_04402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09902__I (.I(_04402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09678__A4 (.I(_04402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09897__A1 (.I(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09730__A1 (.I(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09683__A1 (.I(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10027__A1 (.I(_04404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09748__A1 (.I(_04404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09739__A1 (.I(_04404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09686__A1 (.I(_04404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09682__A1 (.I(_04404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10451__A1 (.I(_04407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10079__A1 (.I(_04407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10075__A1 (.I(_04407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09683__A2 (.I(_04407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10060__A1 (.I(_04411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10012__A2 (.I(_04411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09813__A1 (.I(_04411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09687__A2 (.I(_04411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09827__A1 (.I(_04412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09765__A1 (.I(_04412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09736__A1 (.I(_04412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09797__A1 (.I(_04415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09691__I (.I(_04415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10035__A1 (.I(_04416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09835__A1 (.I(_04416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09790__A1 (.I(_04416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09733__A1 (.I(_04416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09710__A1 (.I(_04416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09807__S (.I(_04417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09702__S (.I(_04417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09701__S (.I(_04417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09695__S (.I(_04417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09693__S (.I(_04417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09797__A2 (.I(_04418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09733__A2 (.I(_04418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09719__A2 (.I(_04418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09713__A2 (.I(_04418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09694__I (.I(_04418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10470__A1 (.I(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10030__C (.I(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09954__A1 (.I(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09853__B2 (.I(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09710__A2 (.I(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10076__A1 (.I(_04420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09981__A1 (.I(_04420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09950__B2 (.I(_04420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09868__A1 (.I(_04420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09696__I (.I(_04420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09820__A1 (.I(_04421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09793__I (.I(_04421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09704__A1 (.I(_04421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09938__B (.I(_04423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09820__A2 (.I(_04423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09801__A2 (.I(_04423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09790__B2 (.I(_04423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09704__A2 (.I(_04423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09979__A1 (.I(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09846__A1 (.I(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09744__I (.I(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09703__A1 (.I(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09866__A1 (.I(_04426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09774__I (.I(_04426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09703__A2 (.I(_04426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09960__B (.I(_04427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09830__A1 (.I(_04427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09827__B2 (.I(_04427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09711__I (.I(_04427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09703__A3 (.I(_04427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10060__A2 (.I(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09764__A1 (.I(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09709__A1 (.I(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09802__A1 (.I(_04431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09751__I (.I(_04431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09708__A1 (.I(_04431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09903__A2 (.I(_04432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09851__A1 (.I(_04432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09767__I (.I(_04432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09708__A2 (.I(_04432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10465__A2 (.I(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10029__A3 (.I(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09827__A2 (.I(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09710__A3 (.I(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10036__A1 (.I(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09915__A1 (.I(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09837__A1 (.I(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09804__A1 (.I(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09723__A1 (.I(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09746__I (.I(_04437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09719__A1 (.I(_04437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09713__A1 (.I(_04437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09766__I (.I(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09728__A1 (.I(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09726__A1 (.I(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09718__A1 (.I(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09728__A2 (.I(_04441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09717__I (.I(_04441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10088__B1 (.I(_04443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09951__I (.I(_04443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09907__A1 (.I(_04443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09868__B1 (.I(_04443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09720__A1 (.I(_04443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09829__I (.I(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09731__A1 (.I(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09726__A2 (.I(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10470__A2 (.I(_04452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10016__A2 (.I(_04452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09992__A2 (.I(_04452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09950__A2 (.I(_04452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09735__A1 (.I(_04452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10477__A2 (.I(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09898__A2 (.I(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09827__B1 (.I(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09731__A2 (.I(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09896__I (.I(_04454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09730__A2 (.I(_04454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10065__A2 (.I(_04456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09937__A2 (.I(_04456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09847__A2 (.I(_04456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09833__A2 (.I(_04456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09732__I (.I(_04456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09822__A2 (.I(_04457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09816__A2 (.I(_04457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09804__A2 (.I(_04457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09785__B (.I(_04457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09735__A2 (.I(_04457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09863__A1 (.I(_04458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09734__I (.I(_04458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10111__B2 (.I(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10100__C (.I(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09913__B (.I(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09786__A1 (.I(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09735__B (.I(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09736__C (.I(_04460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09738__B (.I(_04462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10475__S (.I(_04466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10082__C (.I(_04466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10039__B (.I(_04466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09945__C (.I(_04466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09743__I (.I(_04466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11120__A2 (.I(_04467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10571__A2 (.I(_04467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10120__A1 (.I(_04467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10041__B2 (.I(_04467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09760__A1 (.I(_04467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10452__A1 (.I(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09983__A1 (.I(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09854__B2 (.I(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09816__A1 (.I(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09756__A1 (.I(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10451__B2 (.I(_04469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10102__A1 (.I(_04469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10082__A1 (.I(_04469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09945__A1 (.I(_04469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09756__A2 (.I(_04469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09915__C (.I(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09835__A2 (.I(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09763__I (.I(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09749__A2 (.I(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10075__B (.I(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10066__C (.I(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10058__B (.I(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10034__C (.I(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09755__A1 (.I(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09852__A1 (.I(_04475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09849__A1 (.I(_04475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09799__A1 (.I(_04475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09762__I (.I(_04475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09754__A1 (.I(_04475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09780__A2 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09753__I (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10014__A1 (.I(_04477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09851__A2 (.I(_04477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09818__A2 (.I(_04477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09804__C2 (.I(_04477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09754__A2 (.I(_04477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09809__A2 (.I(_04479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09756__B (.I(_04479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09760__A2 (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10456__B2 (.I(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10056__A3 (.I(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09791__A2 (.I(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09778__A2 (.I(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09759__A2 (.I(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09963__A2 (.I(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09916__A1 (.I(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09817__A1 (.I(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09773__A1 (.I(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09772__A1 (.I(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09958__A2 (.I(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09917__A1 (.I(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09823__A1 (.I(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09817__A2 (.I(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09773__A2 (.I(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09983__C (.I(_04486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09963__B1 (.I(_04486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09854__A1 (.I(_04486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09827__C (.I(_04486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09765__A2 (.I(_04486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10478__B (.I(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10028__A1 (.I(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09765__A3 (.I(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10032__A2 (.I(_04489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09940__I (.I(_04489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09905__A2 (.I(_04489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09903__A1 (.I(_04489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09768__A1 (.I(_04489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10069__A1 (.I(_04490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10060__A3 (.I(_04490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09941__A2 (.I(_04490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09849__A2 (.I(_04490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09768__A2 (.I(_04490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10479__A2 (.I(_04491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10459__B1 (.I(_04491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10028__A2 (.I(_04491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09830__A3 (.I(_04491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09769__A2 (.I(_04491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10461__A1 (.I(_04492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09981__A2 (.I(_04492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09960__A1 (.I(_04492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09785__C (.I(_04492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09772__A2 (.I(_04492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10479__A1 (.I(_04493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09818__A1 (.I(_04493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09817__C (.I(_04493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09775__A2 (.I(_04493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09771__A2 (.I(_04493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11121__A1 (.I(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10463__A1 (.I(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09997__A1 (.I(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09986__A1 (.I(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09772__B (.I(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09795__A2 (.I(_04495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09773__C (.I(_04495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09779__A1 (.I(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10458__A1 (.I(_04497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09991__A1 (.I(_04497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09865__A1 (.I(_04497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09822__A1 (.I(_04497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09778__B1 (.I(_04497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10456__A2 (.I(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10010__A1 (.I(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10000__A1 (.I(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09795__B1 (.I(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09778__B2 (.I(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10077__A2 (.I(_04502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10033__A2 (.I(_04502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09937__B1 (.I(_04502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09814__A2 (.I(_04502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09781__I (.I(_04502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10448__A2 (.I(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10013__C (.I(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09822__B1 (.I(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09804__B1 (.I(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09785__A1 (.I(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10012__A1 (.I(_04505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10005__I (.I(_04505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09941__A1 (.I(_04505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09815__A1 (.I(_04505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09784__A2 (.I(_04505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09791__B1 (.I(_04508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10458__A2 (.I(_04509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10059__A1 (.I(_04509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10033__B2 (.I(_04509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09868__A2 (.I(_04509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09788__I (.I(_04509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10471__A1 (.I(_04510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10452__A2 (.I(_04510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10036__A2 (.I(_04510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09953__A2 (.I(_04510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09790__A2 (.I(_04510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11310__A1 (.I(_04511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10113__A1 (.I(_04511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10102__C (.I(_04511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10093__C (.I(_04511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09790__C (.I(_04511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10459__B2 (.I(_04514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09954__A2 (.I(_04514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09815__A2 (.I(_04514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09801__A1 (.I(_04514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09795__B2 (.I(_04514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10480__A1 (.I(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10468__B2 (.I(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09971__A2 (.I(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09824__A1 (.I(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09811__A1 (.I(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10465__A1 (.I(_04518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10451__A2 (.I(_04518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10079__A2 (.I(_04518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09864__A1 (.I(_04518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09810__A1 (.I(_04518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10460__A2 (.I(_04520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09996__A3 (.I(_04520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09942__C (.I(_04520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09917__C1 (.I(_04520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09810__A2 (.I(_04520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09804__B2 (.I(_04521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09992__B1 (.I(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09983__B1 (.I(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09915__B1 (.I(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09837__A2 (.I(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09804__C1 (.I(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10472__A1 (.I(_04525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09861__A1 (.I(_04525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09823__B1 (.I(_04525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09817__B1 (.I(_04525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09810__B2 (.I(_04525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10109__B (.I(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10067__C (.I(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09944__C (.I(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09870__A2 (.I(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09809__A1 (.I(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09908__A2 (.I(_04527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09905__A1 (.I(_04527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09847__A1 (.I(_04527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09832__I (.I(_04527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09808__I (.I(_04527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09992__B2 (.I(_04528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09963__A1 (.I(_04528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09961__A1 (.I(_04528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09913__A1 (.I(_04528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09809__B (.I(_04528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10051__B2 (.I(_04531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09812__B (.I(_04531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10117__A1 (.I(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10064__A1 (.I(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09822__C (.I(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09816__B (.I(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09817__B2 (.I(_04535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10054__B2 (.I(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09819__B (.I(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09823__B2 (.I(_04540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10057__A1 (.I(_04542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09825__B (.I(_04542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10477__A1 (.I(_04545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09980__A1 (.I(_04545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09962__A1 (.I(_04545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09848__A1 (.I(_04545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09834__A1 (.I(_04545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09959__A1 (.I(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09907__A2 (.I(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09904__A1 (.I(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09898__A1 (.I(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09830__A2 (.I(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10099__A1 (.I(_04548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10059__A2 (.I(_04548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10006__A2 (.I(_04548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09912__A2 (.I(_04548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09833__A1 (.I(_04548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10031__A1 (.I(_04549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10029__A2 (.I(_04549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09937__A1 (.I(_04549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09899__A1 (.I(_04549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09833__B (.I(_04549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10107__A1 (.I(_04550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10099__B (.I(_04550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10090__A1 (.I(_04550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09834__A3 (.I(_04550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09839__A2 (.I(_04551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10088__C (.I(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10074__B (.I(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10063__A1 (.I(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09943__B (.I(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09837__B (.I(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10008__C (.I(_04555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09839__A4 (.I(_04555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09840__B (.I(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10048__B2 (.I(_04557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09928__C (.I(_04557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09841__B (.I(_04557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10119__B1 (.I(_04558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09987__C2 (.I(_04558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09956__C2 (.I(_04558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09871__A1 (.I(_04558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09857__A1 (.I(_04558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09857__A2 (.I(_04559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10471__A2 (.I(_04560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10453__A1 (.I(_04560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10450__B (.I(_04560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09954__B1 (.I(_04560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09855__A1 (.I(_04560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10077__A1 (.I(_04561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10031__A2 (.I(_04561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09912__B1 (.I(_04561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09866__A2 (.I(_04561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09846__A2 (.I(_04561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10449__A1 (.I(_04562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09855__A2 (.I(_04562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09978__A1 (.I(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09962__A2 (.I(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09862__A1 (.I(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09861__A2 (.I(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09848__A2 (.I(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10448__A1 (.I(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09983__A2 (.I(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09979__A2 (.I(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09915__A2 (.I(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09853__A2 (.I(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10478__A1 (.I(_04567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09961__A2 (.I(_04567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09910__A1 (.I(_04567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09852__A2 (.I(_04567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09862__A2 (.I(_04568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09853__B1 (.I(_04568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09857__B1 (.I(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10094__A2 (.I(_04572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10083__A2 (.I(_04572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10069__C (.I(_04572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09946__A2 (.I(_04572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09857__B2 (.I(_04572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09931__A1 (.I(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09858__B (.I(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09871__A2 (.I(_04574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09868__B2 (.I(_04574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10478__C (.I(_04575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10092__C (.I(_04575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09996__A2 (.I(_04575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09985__C (.I(_04575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09869__A1 (.I(_04575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09869__A2 (.I(_04580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10461__C (.I(_04581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09869__B1 (.I(_04581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10470__C (.I(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10036__C (.I(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10003__A2 (.I(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09944__A1 (.I(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09868__C (.I(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10038__B2 (.I(_04585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09964__A1 (.I(_04585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09955__A1 (.I(_04585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09919__C (.I(_04585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09871__B2 (.I(_04585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09935__B2 (.I(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09872__B (.I(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09917__B2 (.I(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09894__A2 (.I(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10065__A1 (.I(_04601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09943__A1 (.I(_04601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09917__A2 (.I(_04601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09912__B2 (.I(_04601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09901__A1 (.I(_04601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10448__B (.I(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10077__B (.I(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10074__A1 (.I(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09982__I (.I(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09897__A2 (.I(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10038__A1 (.I(_04608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10036__B2 (.I(_04608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09917__C2 (.I(_04608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09915__B2 (.I(_04608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09912__A1 (.I(_04608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10074__C (.I(_04609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10063__A2 (.I(_04609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09985__A2 (.I(_04609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09943__A2 (.I(_04609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09904__A2 (.I(_04609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10117__A3 (.I(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10006__B (.I(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09961__B (.I(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09910__B (.I(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10120__A2 (.I(_04619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10017__B (.I(_04619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10007__B (.I(_04619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09993__B (.I(_04619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09914__B (.I(_04619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09919__A1 (.I(_04620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09920__A2 (.I(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09977__A1 (.I(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09921__B (.I(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09934__A2 (.I(_04627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09929__A2 (.I(_04627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09923__A2 (.I(_04627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09948__A1 (.I(_04629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09947__A2 (.I(_04629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09935__A2 (.I(_04629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09930__A2 (.I(_04629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09928__A1 (.I(_04629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10481__A2 (.I(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10464__A2 (.I(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10119__A2 (.I(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10070__A2 (.I(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09926__A2 (.I(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10446__A2 (.I(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10053__A2 (.I(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10050__A2 (.I(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10047__A2 (.I(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09934__B (.I(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09944__A2 (.I(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09948__A2 (.I(_04647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10480__A2 (.I(_04650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10111__A1 (.I(_04650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10106__A1 (.I(_04650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09953__A1 (.I(_04650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09950__A1 (.I(_04650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09957__A1 (.I(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10452__B1 (.I(_04652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10073__A1 (.I(_04652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10036__B1 (.I(_04652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09985__B2 (.I(_04652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09953__B1 (.I(_04652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09956__C1 (.I(_04653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09953__B2 (.I(_04653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09957__B (.I(_04657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09979__A3 (.I(_04659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09960__A2 (.I(_04659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09963__C (.I(_04662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09964__A2 (.I(_04663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09998__A3 (.I(_04665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09966__A2 (.I(_04665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10009__A2 (.I(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09999__A2 (.I(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09971__B (.I(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10019__A2 (.I(_04672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09987__A2 (.I(_04672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09976__A2 (.I(_04672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09973__A2 (.I(_04672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09986__A2 (.I(_04679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10456__A1 (.I(_04680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10452__B2 (.I(_04680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10016__A1 (.I(_04680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09985__A1 (.I(_04680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09983__B2 (.I(_04680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09986__A3 (.I(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09987__C1 (.I(_04682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09985__B1 (.I(_04682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09988__A1 (.I(_04684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09997__A2 (.I(_04690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10467__A1 (.I(_04692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10459__A1 (.I(_04692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10092__A1 (.I(_04692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10058__A1 (.I(_04692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09996__A1 (.I(_04692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10000__B (.I(_04694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10461__B (.I(_04700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10449__A2 (.I(_04700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10100__A2 (.I(_04700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10090__A2 (.I(_04700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10007__A1 (.I(_04700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10471__B2 (.I(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10100__A1 (.I(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10098__A1 (.I(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10013__A2 (.I(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10006__A1 (.I(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10008__B (.I(_04703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10010__B (.I(_04704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10117__A2 (.I(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10106__A2 (.I(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10066__A2 (.I(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10034__A2 (.I(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10016__B (.I(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10018__B1 (.I(_04712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10572__A1 (.I(_04713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10025__A1 (.I(_04713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10048__A1 (.I(_04715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10023__A1 (.I(_04715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10068__A1 (.I(_04721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10066__A1 (.I(_04721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10034__A1 (.I(_04721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10032__A1 (.I(_04721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10030__A1 (.I(_04721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10035__B (.I(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10037__A1 (.I(_04729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10447__B2 (.I(_04732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10041__A1 (.I(_04732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10056__A4 (.I(_04736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10044__A2 (.I(_04736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10084__I (.I(_04737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10053__B (.I(_04737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10050__B (.I(_04737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10046__I (.I(_04737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10045__I (.I(_04737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10086__A1 (.I(_04738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10071__A2 (.I(_04738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10054__A2 (.I(_04738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10051__A2 (.I(_04738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10048__A2 (.I(_04738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10115__A2 (.I(_04739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10104__A2 (.I(_04739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10070__B (.I(_04739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10055__A2 (.I(_04739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10047__B (.I(_04739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10057__A3 (.I(_04746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10111__A2 (.I(_04750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10098__A2 (.I(_04750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10062__B (.I(_04750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10069__B (.I(_04757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10082__A2 (.I(_04760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10073__A2 (.I(_04760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10080__B (.I(_04767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10081__C (.I(_04768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10093__B2 (.I(_04779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10096__A2 (.I(_04780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10101__A2 (.I(_04786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10105__A2 (.I(_04788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10111__C (.I(_04795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10116__A2 (.I(_04796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10116__A3 (.I(_04799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10120__A3 (.I(_04801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10850__I (.I(_04807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10741__I (.I(_04807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10632__I (.I(_04807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10483__I (.I(_04807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10126__I (.I(_04807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10427__A1 (.I(_04808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10371__A1 (.I(_04808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10264__A1 (.I(_04808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10165__A1 (.I(_04808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10131__A1 (.I(_04808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10159__A2 (.I(_04809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10138__I (.I(_04809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10129__I (.I(_04809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10128__I (.I(_04809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10160__A2 (.I(_04811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10156__A2 (.I(_04811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10152__A2 (.I(_04811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10134__A2 (.I(_04811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10130__A2 (.I(_04811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10856__I (.I(_04813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10747__I (.I(_04813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10638__I (.I(_04813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10489__I (.I(_04813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10133__I (.I(_04813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10429__A1 (.I(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10373__A1 (.I(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10266__A1 (.I(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10167__A1 (.I(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10135__A1 (.I(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10859__I (.I(_04816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10750__I (.I(_04816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10641__I (.I(_04816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10492__I (.I(_04816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10137__I (.I(_04816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10432__A1 (.I(_04817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10376__A1 (.I(_04817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10269__A1 (.I(_04817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10170__A1 (.I(_04817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10140__A1 (.I(_04817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10434__A1 (.I(_04821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10378__A1 (.I(_04821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10271__A1 (.I(_04821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10172__A1 (.I(_04821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10144__A1 (.I(_04821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10436__A1 (.I(_04824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10380__A1 (.I(_04824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10273__A1 (.I(_04824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10174__A1 (.I(_04824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10148__A1 (.I(_04824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10869__I (.I(_04826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10760__I (.I(_04826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10651__I (.I(_04826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10502__I (.I(_04826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10150__I (.I(_04826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10438__A1 (.I(_04827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10382__A1 (.I(_04827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10275__A1 (.I(_04827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10176__A1 (.I(_04827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10152__A1 (.I(_04827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10872__I (.I(_04829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10763__I (.I(_04829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10654__I (.I(_04829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10505__I (.I(_04829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10154__I (.I(_04829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10440__A1 (.I(_04830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10384__A1 (.I(_04830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10277__A1 (.I(_04830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10178__A1 (.I(_04830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10156__A1 (.I(_04830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10875__I (.I(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10766__I (.I(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10657__I (.I(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10508__I (.I(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10158__I (.I(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10442__A1 (.I(_04833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10386__A1 (.I(_04833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10279__A1 (.I(_04833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10180__A1 (.I(_04833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10160__A1 (.I(_04833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10174__A2 (.I(_04836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10172__A2 (.I(_04836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10170__A2 (.I(_04836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10167__A2 (.I(_04836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10165__A2 (.I(_04836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10180__A2 (.I(_04837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10178__A2 (.I(_04837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10176__A2 (.I(_04837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10166__A2 (.I(_04837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10164__A2 (.I(_04837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10177__A2 (.I(_04840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10175__A2 (.I(_04840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10173__A2 (.I(_04840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10171__A2 (.I(_04840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10169__A2 (.I(_04840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10243__S (.I(_04848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10241__S (.I(_04848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10239__S (.I(_04848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10195__I (.I(_04848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10184__I (.I(_04848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10193__S (.I(_04849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10191__S (.I(_04849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10189__S (.I(_04849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10187__S (.I(_04849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10185__S (.I(_04849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10204__S (.I(_04855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10202__S (.I(_04855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10200__S (.I(_04855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10198__S (.I(_04855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10196__S (.I(_04855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10215__S (.I(_04861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10213__S (.I(_04861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10211__S (.I(_04861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10209__S (.I(_04861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10207__S (.I(_04861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10226__S (.I(_04867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10224__S (.I(_04867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10222__S (.I(_04867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10220__S (.I(_04867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10218__S (.I(_04867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10257__A1 (.I(_04886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10251__B1 (.I(_04886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10259__A2 (.I(_04888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10258__A1 (.I(_04888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10255__A2 (.I(_04888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10254__A2 (.I(_04888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10278__A2 (.I(_04893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10267__I (.I(_04893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10262__I (.I(_04893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10261__I (.I(_04893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10273__A2 (.I(_04894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10271__A2 (.I(_04894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10269__A2 (.I(_04894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10266__A2 (.I(_04894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10264__A2 (.I(_04894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10279__A2 (.I(_04895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10277__A2 (.I(_04895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10275__A2 (.I(_04895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10265__A2 (.I(_04895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10263__A2 (.I(_04895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10276__A2 (.I(_04898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10274__A2 (.I(_04898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10272__A2 (.I(_04898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10270__A2 (.I(_04898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10268__A2 (.I(_04898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10342__I (.I(_04905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10330__I (.I(_04905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10318__I (.I(_04905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10306__I (.I(_04905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10281__I (.I(_04905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10363__A2 (.I(_04906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10356__A2 (.I(_04906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10354__A2 (.I(_04906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10294__I (.I(_04906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10282__I (.I(_04906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11312__A1 (.I(_04907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10292__A2 (.I(_04907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10290__A2 (.I(_04907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10288__A2 (.I(_04907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10286__A2 (.I(_04907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10345__I (.I(_04908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10333__I (.I(_04908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10321__I (.I(_04908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10284__I (.I(_04908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10363__B1 (.I(_04909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10356__B1 (.I(_04909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10309__I (.I(_04909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10297__I (.I(_04909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10285__I (.I(_04909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10295__B1 (.I(_04910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10292__B1 (.I(_04910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10290__B1 (.I(_04910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10288__B1 (.I(_04910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10286__B1 (.I(_04910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10304__A2 (.I(_04915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10302__A2 (.I(_04915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10300__A2 (.I(_04915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10298__A2 (.I(_04915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10295__A2 (.I(_04915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10328__A2 (.I(_04929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10326__A2 (.I(_04929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10324__A2 (.I(_04929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10322__A2 (.I(_04929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10319__A2 (.I(_04929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10331__B1 (.I(_04931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10328__B1 (.I(_04931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10326__B1 (.I(_04931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10324__B1 (.I(_04931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10322__B1 (.I(_04931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10340__A2 (.I(_04936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10338__A2 (.I(_04936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10336__A2 (.I(_04936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10334__A2 (.I(_04936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10331__A2 (.I(_04936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10343__B1 (.I(_04938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10340__B1 (.I(_04938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10338__B1 (.I(_04938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10336__B1 (.I(_04938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10334__B1 (.I(_04938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10354__B1 (.I(_04945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10352__B1 (.I(_04945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10350__B1 (.I(_04945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10348__B1 (.I(_04945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10346__B1 (.I(_04945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11117__A1 (.I(_04952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11115__A1 (.I(_04952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10359__A1 (.I(_04952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10362__A1 (.I(_04953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10361__B (.I(_04953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10363__B2 (.I(_04956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11250__A2 (.I(_04958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10809__I (.I(_04958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10680__I (.I(_04958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10366__I (.I(_04958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10380__A2 (.I(_04961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10378__A2 (.I(_04961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10376__A2 (.I(_04961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10373__A2 (.I(_04961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10371__A2 (.I(_04961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10386__A2 (.I(_04962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10384__A2 (.I(_04962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10382__A2 (.I(_04962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10372__A2 (.I(_04962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10370__A2 (.I(_04962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10383__A2 (.I(_04965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10381__A2 (.I(_04965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10379__A2 (.I(_04965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10377__A2 (.I(_04965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10375__A2 (.I(_04965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10403__S (.I(_04972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10401__S (.I(_04972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10399__S (.I(_04972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10388__I (.I(_04972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10397__S (.I(_04973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10395__S (.I(_04973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10393__S (.I(_04973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10391__S (.I(_04973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10389__S (.I(_04973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10421__S (.I(_04982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10419__S (.I(_04982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10417__S (.I(_04982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10406__I (.I(_04982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10415__S (.I(_04983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10413__S (.I(_04983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10411__S (.I(_04983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10409__S (.I(_04983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10407__S (.I(_04983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10441__A2 (.I(_04992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10430__I (.I(_04992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10425__I (.I(_04992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10424__I (.I(_04992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10436__A2 (.I(_04993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10434__A2 (.I(_04993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10432__A2 (.I(_04993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10429__A2 (.I(_04993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10427__A2 (.I(_04993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10474__A2 (.I(_05004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10473__A2 (.I(_05004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10455__S (.I(_05004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10444__A2 (.I(_05004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10451__B1 (.I(_05010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10454__A2 (.I(_05011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10464__B (.I(_05022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10470__B (.I(_05025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10467__A2 (.I(_05025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10475__I0 (.I(_05030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10482__B1 (.I(_05037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10581__A1 (.I(_05039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10555__A1 (.I(_05039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10535__A1 (.I(_05039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10515__A1 (.I(_05039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10488__A1 (.I(_05039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10509__A2 (.I(_05040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10493__I (.I(_05040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10486__I (.I(_05040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10485__I (.I(_05040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10510__A2 (.I(_05042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10507__A2 (.I(_05042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10504__A2 (.I(_05042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10490__A2 (.I(_05042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10487__A2 (.I(_05042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10583__A1 (.I(_05044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10557__A1 (.I(_05044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10537__A1 (.I(_05044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10517__A1 (.I(_05044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10491__A1 (.I(_05044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10586__A1 (.I(_05046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10560__A1 (.I(_05046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10540__A1 (.I(_05046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10520__A1 (.I(_05046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10495__A1 (.I(_05046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10506__A2 (.I(_05047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10503__A2 (.I(_05047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10500__A2 (.I(_05047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10497__A2 (.I(_05047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10494__A2 (.I(_05047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10588__A1 (.I(_05049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10562__A1 (.I(_05049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10542__A1 (.I(_05049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10522__A1 (.I(_05049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10498__A1 (.I(_05049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10590__A1 (.I(_05051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10564__A1 (.I(_05051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10544__A1 (.I(_05051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10524__A1 (.I(_05051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10501__A1 (.I(_05051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10592__A1 (.I(_05053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10566__A1 (.I(_05053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10546__A1 (.I(_05053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10526__A1 (.I(_05053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10504__A1 (.I(_05053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10594__A1 (.I(_05055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10568__A1 (.I(_05055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10548__A1 (.I(_05055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10528__A1 (.I(_05055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10507__A1 (.I(_05055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10596__A1 (.I(_05057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10570__A1 (.I(_05057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10550__A1 (.I(_05057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10530__A1 (.I(_05057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10510__A1 (.I(_05057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10529__A2 (.I(_05059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10518__I (.I(_05059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10513__I (.I(_05059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10512__I (.I(_05059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10524__A2 (.I(_05060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10522__A2 (.I(_05060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10520__A2 (.I(_05060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10517__A2 (.I(_05060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10515__A2 (.I(_05060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10527__A2 (.I(_05064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10525__A2 (.I(_05064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10523__A2 (.I(_05064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10521__A2 (.I(_05064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10519__A2 (.I(_05064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10549__A2 (.I(_05071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10538__I (.I(_05071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10533__I (.I(_05071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10532__I (.I(_05071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10544__A2 (.I(_05072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10542__A2 (.I(_05072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10540__A2 (.I(_05072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10537__A2 (.I(_05072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10535__A2 (.I(_05072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10550__A2 (.I(_05073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10548__A2 (.I(_05073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10546__A2 (.I(_05073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10536__A2 (.I(_05073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10534__A2 (.I(_05073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10547__A2 (.I(_05076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10545__A2 (.I(_05076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10543__A2 (.I(_05076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10541__A2 (.I(_05076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10539__A2 (.I(_05076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10569__A2 (.I(_05083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10558__I (.I(_05083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10553__I (.I(_05083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10552__I (.I(_05083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10567__A2 (.I(_05088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10565__A2 (.I(_05088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10563__A2 (.I(_05088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10561__A2 (.I(_05088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10559__A2 (.I(_05088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11192__A1 (.I(_05098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11172__A1 (.I(_05098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11152__A1 (.I(_05098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11125__A1 (.I(_05098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10577__A1 (.I(_05098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10595__A2 (.I(_05099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10584__I (.I(_05099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10579__I (.I(_05099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10578__I (.I(_05099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10593__A2 (.I(_05104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10591__A2 (.I(_05104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10589__A2 (.I(_05104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10587__A2 (.I(_05104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10585__A2 (.I(_05104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10606__S (.I(_05111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10604__S (.I(_05111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10602__S (.I(_05111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10600__S (.I(_05111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10598__S (.I(_05111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10617__S (.I(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10615__S (.I(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10613__S (.I(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10611__S (.I(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10609__S (.I(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10725__A1 (.I(_05130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10705__A1 (.I(_05130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10685__A1 (.I(_05130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10664__A1 (.I(_05130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10637__A1 (.I(_05130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10658__A2 (.I(_05131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10642__I (.I(_05131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10635__I (.I(_05131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10634__I (.I(_05131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10650__A2 (.I(_05132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10647__A2 (.I(_05132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10644__A2 (.I(_05132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10640__A2 (.I(_05132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10637__A2 (.I(_05132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10659__A2 (.I(_05133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10656__A2 (.I(_05133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10653__A2 (.I(_05133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10639__A2 (.I(_05133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10636__A2 (.I(_05133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10727__A1 (.I(_05135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10707__A1 (.I(_05135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10687__A1 (.I(_05135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10666__A1 (.I(_05135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10640__A1 (.I(_05135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10730__A1 (.I(_05137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10710__A1 (.I(_05137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10690__A1 (.I(_05137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10669__A1 (.I(_05137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10644__A1 (.I(_05137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10655__A2 (.I(_05138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10652__A2 (.I(_05138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10649__A2 (.I(_05138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10646__A2 (.I(_05138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10643__A2 (.I(_05138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10732__A1 (.I(_05140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10712__A1 (.I(_05140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10692__A1 (.I(_05140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10671__A1 (.I(_05140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10647__A1 (.I(_05140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10734__A1 (.I(_05142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10714__A1 (.I(_05142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10694__A1 (.I(_05142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10673__A1 (.I(_05142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10650__A1 (.I(_05142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10736__A1 (.I(_05144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10716__A1 (.I(_05144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10696__A1 (.I(_05144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10675__A1 (.I(_05144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10653__A1 (.I(_05144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10738__A1 (.I(_05146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10718__A1 (.I(_05146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10698__A1 (.I(_05146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10677__A1 (.I(_05146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10656__A1 (.I(_05146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10740__A1 (.I(_05148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10720__A1 (.I(_05148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10700__A1 (.I(_05148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10679__A1 (.I(_05148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10659__A1 (.I(_05148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10678__A2 (.I(_05150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10667__I (.I(_05150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10662__I (.I(_05150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10661__I (.I(_05150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10673__A2 (.I(_05151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10671__A2 (.I(_05151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10669__A2 (.I(_05151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10666__A2 (.I(_05151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10664__A2 (.I(_05151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10679__A2 (.I(_05152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10677__A2 (.I(_05152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10675__A2 (.I(_05152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10665__A2 (.I(_05152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10663__A2 (.I(_05152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10789__A2 (.I(_05162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10769__A2 (.I(_05162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10721__A2 (.I(_05162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10701__A2 (.I(_05162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10681__A2 (.I(_05162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10699__A2 (.I(_05163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10688__I (.I(_05163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10683__I (.I(_05163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10682__I (.I(_05163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10700__A2 (.I(_05165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10698__A2 (.I(_05165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10696__A2 (.I(_05165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10686__A2 (.I(_05165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10684__A2 (.I(_05165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10697__A2 (.I(_05168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10695__A2 (.I(_05168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10693__A2 (.I(_05168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10691__A2 (.I(_05168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10689__A2 (.I(_05168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10719__A2 (.I(_05175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10708__I (.I(_05175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10703__I (.I(_05175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10702__I (.I(_05175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10714__A2 (.I(_05176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10712__A2 (.I(_05176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10710__A2 (.I(_05176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10707__A2 (.I(_05176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10705__A2 (.I(_05176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10720__A2 (.I(_05177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10718__A2 (.I(_05177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10716__A2 (.I(_05177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10706__A2 (.I(_05177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10704__A2 (.I(_05177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10834__A1 (.I(_05199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10814__A1 (.I(_05199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10793__A1 (.I(_05199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10773__A1 (.I(_05199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10746__A1 (.I(_05199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10759__A2 (.I(_05201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10756__A2 (.I(_05201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10753__A2 (.I(_05201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10749__A2 (.I(_05201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10746__A2 (.I(_05201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10836__A1 (.I(_05204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10816__A1 (.I(_05204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10795__A1 (.I(_05204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10775__A1 (.I(_05204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10749__A1 (.I(_05204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10839__A1 (.I(_05206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10819__A1 (.I(_05206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10798__A1 (.I(_05206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10778__A1 (.I(_05206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10753__A1 (.I(_05206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10764__A2 (.I(_05207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10761__A2 (.I(_05207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10758__A2 (.I(_05207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10755__A2 (.I(_05207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10752__A2 (.I(_05207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10841__A1 (.I(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10821__A1 (.I(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10800__A1 (.I(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10780__A1 (.I(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10756__A1 (.I(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10843__A1 (.I(_05211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10823__A1 (.I(_05211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10802__A1 (.I(_05211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10782__A1 (.I(_05211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10759__A1 (.I(_05211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10845__A1 (.I(_05213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10825__A1 (.I(_05213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10804__A1 (.I(_05213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10784__A1 (.I(_05213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10762__A1 (.I(_05213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10847__A1 (.I(_05215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10827__A1 (.I(_05215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10806__A1 (.I(_05215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10786__A1 (.I(_05215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10765__A1 (.I(_05215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10849__A1 (.I(_05217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10829__A1 (.I(_05217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10808__A1 (.I(_05217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10788__A1 (.I(_05217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10768__A1 (.I(_05217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10787__A2 (.I(_05219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10776__I (.I(_05219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10771__I (.I(_05219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10770__I (.I(_05219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10782__A2 (.I(_05220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10780__A2 (.I(_05220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10778__A2 (.I(_05220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10775__A2 (.I(_05220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10773__A2 (.I(_05220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10788__A2 (.I(_05221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10786__A2 (.I(_05221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10784__A2 (.I(_05221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10774__A2 (.I(_05221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10772__A2 (.I(_05221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10785__A2 (.I(_05224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10783__A2 (.I(_05224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10781__A2 (.I(_05224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10779__A2 (.I(_05224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10777__A2 (.I(_05224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10807__A2 (.I(_05231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10796__I (.I(_05231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10791__I (.I(_05231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10790__I (.I(_05231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10802__A2 (.I(_05232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10800__A2 (.I(_05232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10798__A2 (.I(_05232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10795__A2 (.I(_05232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10793__A2 (.I(_05232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10808__A2 (.I(_05233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10806__A2 (.I(_05233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10804__A2 (.I(_05233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10794__A2 (.I(_05233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10792__A2 (.I(_05233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10805__A2 (.I(_05236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10803__A2 (.I(_05236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10801__A2 (.I(_05236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10799__A2 (.I(_05236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10797__A2 (.I(_05236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11230__A2 (.I(_05243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11025__A2 (.I(_05243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10978__A2 (.I(_05243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10851__A2 (.I(_05243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10810__A2 (.I(_05243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10828__A2 (.I(_05244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10817__I (.I(_05244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10812__I (.I(_05244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10811__I (.I(_05244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10823__A2 (.I(_05245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10821__A2 (.I(_05245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10819__A2 (.I(_05245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10816__A2 (.I(_05245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10814__A2 (.I(_05245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10829__A2 (.I(_05246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10827__A2 (.I(_05246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10825__A2 (.I(_05246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10815__A2 (.I(_05246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10813__A2 (.I(_05246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10826__A2 (.I(_05249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10824__A2 (.I(_05249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10822__A2 (.I(_05249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10820__A2 (.I(_05249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10818__A2 (.I(_05249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10843__A2 (.I(_05257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10841__A2 (.I(_05257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10839__A2 (.I(_05257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10836__A2 (.I(_05257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10834__A2 (.I(_05257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10846__A2 (.I(_05261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10844__A2 (.I(_05261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10842__A2 (.I(_05261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10840__A2 (.I(_05261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10838__A2 (.I(_05261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10961__A1 (.I(_05268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10923__A1 (.I(_05268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10903__A1 (.I(_05268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10882__A1 (.I(_05268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10855__A1 (.I(_05268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10868__A2 (.I(_05270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10865__A2 (.I(_05270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10862__A2 (.I(_05270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10858__A2 (.I(_05270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10855__A2 (.I(_05270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10963__A1 (.I(_05273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10925__A1 (.I(_05273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10905__A1 (.I(_05273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10884__A1 (.I(_05273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10858__A1 (.I(_05273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10966__A1 (.I(_05275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10928__A1 (.I(_05275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10908__A1 (.I(_05275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10887__A1 (.I(_05275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10862__A1 (.I(_05275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10873__A2 (.I(_05276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10870__A2 (.I(_05276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10867__A2 (.I(_05276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10864__A2 (.I(_05276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10861__A2 (.I(_05276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10968__A1 (.I(_05278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10930__A1 (.I(_05278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10910__A1 (.I(_05278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10889__A1 (.I(_05278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10865__A1 (.I(_05278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10970__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10932__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10912__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10891__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10868__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10972__A1 (.I(_05282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10934__A1 (.I(_05282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10914__A1 (.I(_05282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10893__A1 (.I(_05282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10871__A1 (.I(_05282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10974__A1 (.I(_05284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10936__A1 (.I(_05284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10916__A1 (.I(_05284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10895__A1 (.I(_05284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10874__A1 (.I(_05284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10976__A1 (.I(_05286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10938__A1 (.I(_05286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10918__A1 (.I(_05286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10897__A1 (.I(_05286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10877__A1 (.I(_05286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10891__A2 (.I(_05289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10889__A2 (.I(_05289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10887__A2 (.I(_05289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10884__A2 (.I(_05289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10882__A2 (.I(_05289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10897__A2 (.I(_05290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10895__A2 (.I(_05290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10893__A2 (.I(_05290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10883__A2 (.I(_05290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10881__A2 (.I(_05290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10894__A2 (.I(_05293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10892__A2 (.I(_05293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10890__A2 (.I(_05293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10888__A2 (.I(_05293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10886__A2 (.I(_05293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11065__A1 (.I(_05300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11045__A1 (.I(_05300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11005__A1 (.I(_05300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10957__A1 (.I(_05300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10899__A1 (.I(_05300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10912__A2 (.I(_05302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10910__A2 (.I(_05302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10908__A2 (.I(_05302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10905__A2 (.I(_05302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10903__A2 (.I(_05302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10918__A2 (.I(_05303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10916__A2 (.I(_05303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10914__A2 (.I(_05303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10904__A2 (.I(_05303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10902__A2 (.I(_05303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10935__A2 (.I(_05318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10933__A2 (.I(_05318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10931__A2 (.I(_05318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10929__A2 (.I(_05318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10927__A2 (.I(_05318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10955__S (.I(_05325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10953__S (.I(_05325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10951__S (.I(_05325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10940__I (.I(_05325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10949__S (.I(_05326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10947__S (.I(_05326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10945__S (.I(_05326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10943__S (.I(_05326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10941__S (.I(_05326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10970__A2 (.I(_05336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10968__A2 (.I(_05336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10966__A2 (.I(_05336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10963__A2 (.I(_05336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10961__A2 (.I(_05336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10976__A2 (.I(_05337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10974__A2 (.I(_05337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10972__A2 (.I(_05337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10962__A2 (.I(_05337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10960__A2 (.I(_05337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10973__A2 (.I(_05340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10971__A2 (.I(_05340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10969__A2 (.I(_05340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10967__A2 (.I(_05340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10965__A2 (.I(_05340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11069__A1 (.I(_05347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11049__A1 (.I(_05347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11029__A1 (.I(_05347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11009__A1 (.I(_05347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10982__A1 (.I(_05347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10995__A2 (.I(_05349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10992__A2 (.I(_05349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10989__A2 (.I(_05349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10985__A2 (.I(_05349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10982__A2 (.I(_05349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11071__A1 (.I(_05352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11051__A1 (.I(_05352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11031__A1 (.I(_05352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11011__A1 (.I(_05352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10985__A1 (.I(_05352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11074__A1 (.I(_05354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11054__A1 (.I(_05354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11034__A1 (.I(_05354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11014__A1 (.I(_05354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10989__A1 (.I(_05354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11076__A1 (.I(_05357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11056__A1 (.I(_05357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11036__A1 (.I(_05357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11016__A1 (.I(_05357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10992__A1 (.I(_05357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11078__A1 (.I(_05359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11058__A1 (.I(_05359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11038__A1 (.I(_05359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11018__A1 (.I(_05359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10995__A1 (.I(_05359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11080__A1 (.I(_05361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11060__A1 (.I(_05361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11040__A1 (.I(_05361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11020__A1 (.I(_05361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10998__A1 (.I(_05361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11082__A1 (.I(_05363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11062__A1 (.I(_05363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11042__A1 (.I(_05363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11022__A1 (.I(_05363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11001__A1 (.I(_05363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11084__A1 (.I(_05365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11064__A1 (.I(_05365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11044__A1 (.I(_05365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11024__A1 (.I(_05365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11004__A1 (.I(_05365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11018__A2 (.I(_05368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11016__A2 (.I(_05368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11014__A2 (.I(_05368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11011__A2 (.I(_05368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11009__A2 (.I(_05368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11024__A2 (.I(_05369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11022__A2 (.I(_05369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11020__A2 (.I(_05369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11010__A2 (.I(_05369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11008__A2 (.I(_05369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11021__A2 (.I(_05372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11019__A2 (.I(_05372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11017__A2 (.I(_05372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11015__A2 (.I(_05372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11013__A2 (.I(_05372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11043__A2 (.I(_05379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11032__I (.I(_05379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11027__I (.I(_05379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11026__I (.I(_05379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11038__A2 (.I(_05380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11036__A2 (.I(_05380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11034__A2 (.I(_05380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11031__A2 (.I(_05380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11029__A2 (.I(_05380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11041__A2 (.I(_05384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11039__A2 (.I(_05384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11037__A2 (.I(_05384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11035__A2 (.I(_05384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11033__A2 (.I(_05384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11058__A2 (.I(_05392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11056__A2 (.I(_05392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11054__A2 (.I(_05392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11051__A2 (.I(_05392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11049__A2 (.I(_05392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11064__A2 (.I(_05393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11062__A2 (.I(_05393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11060__A2 (.I(_05393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11050__A2 (.I(_05393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11048__A2 (.I(_05393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11234__A1 (.I(_05444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11196__A1 (.I(_05444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11176__A1 (.I(_05444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11156__A1 (.I(_05444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11129__A1 (.I(_05444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11150__A2 (.I(_05445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11134__I (.I(_05445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11127__I (.I(_05445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11126__I (.I(_05445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11236__A1 (.I(_05449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11198__A1 (.I(_05449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11178__A1 (.I(_05449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11158__A1 (.I(_05449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11132__A1 (.I(_05449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11239__A1 (.I(_05451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11201__A1 (.I(_05451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11181__A1 (.I(_05451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11161__A1 (.I(_05451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11136__A1 (.I(_05451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11147__A2 (.I(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11144__A2 (.I(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11141__A2 (.I(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11138__A2 (.I(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11135__A2 (.I(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11241__A1 (.I(_05454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11203__A1 (.I(_05454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11183__A1 (.I(_05454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11163__A1 (.I(_05454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11139__A1 (.I(_05454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11243__A1 (.I(_05456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11205__A1 (.I(_05456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11185__A1 (.I(_05456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11165__A1 (.I(_05456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11142__A1 (.I(_05456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11245__A1 (.I(_05458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11207__A1 (.I(_05458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11187__A1 (.I(_05458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11167__A1 (.I(_05458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11145__A1 (.I(_05458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11247__A1 (.I(_05460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11209__A1 (.I(_05460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11189__A1 (.I(_05460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11169__A1 (.I(_05460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11148__A1 (.I(_05460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11249__A1 (.I(_05462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11211__A1 (.I(_05462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11191__A1 (.I(_05462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11171__A1 (.I(_05462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11151__A1 (.I(_05462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11170__A2 (.I(_05464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11159__I (.I(_05464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11154__I (.I(_05464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11153__I (.I(_05464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11171__A2 (.I(_05466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11169__A2 (.I(_05466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11167__A2 (.I(_05466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11157__A2 (.I(_05466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11155__A2 (.I(_05466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11168__A2 (.I(_05469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11166__A2 (.I(_05469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11164__A2 (.I(_05469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11162__A2 (.I(_05469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11160__A2 (.I(_05469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11190__A2 (.I(_05476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11179__I (.I(_05476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11174__I (.I(_05476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11173__I (.I(_05476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11185__A2 (.I(_05477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11183__A2 (.I(_05477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11181__A2 (.I(_05477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11178__A2 (.I(_05477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11176__A2 (.I(_05477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11191__A2 (.I(_05478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11189__A2 (.I(_05478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11187__A2 (.I(_05478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11177__A2 (.I(_05478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11175__A2 (.I(_05478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11188__A2 (.I(_05481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11186__A2 (.I(_05481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11184__A2 (.I(_05481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11182__A2 (.I(_05481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11180__A2 (.I(_05481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11208__A2 (.I(_05493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11206__A2 (.I(_05493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11204__A2 (.I(_05493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11202__A2 (.I(_05493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11200__A2 (.I(_05493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11228__S (.I(_05500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11226__S (.I(_05500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11224__S (.I(_05500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11213__I (.I(_05500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11222__S (.I(_05501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11220__S (.I(_05501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11218__S (.I(_05501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11216__S (.I(_05501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11214__S (.I(_05501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11243__A2 (.I(_05511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11241__A2 (.I(_05511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11239__A2 (.I(_05511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11236__A2 (.I(_05511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11234__A2 (.I(_05511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11249__A2 (.I(_05512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11247__A2 (.I(_05512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11245__A2 (.I(_05512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11235__A2 (.I(_05512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11233__A2 (.I(_05512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11246__A2 (.I(_05515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11244__A2 (.I(_05515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11242__A2 (.I(_05515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11240__A2 (.I(_05515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11238__A2 (.I(_05515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11268__A2 (.I(_05522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11257__I (.I(_05522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11252__I (.I(_05522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11251__I (.I(_05522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11263__A2 (.I(_05523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11261__A2 (.I(_05523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11259__A2 (.I(_05523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11256__A2 (.I(_05523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11254__A2 (.I(_05523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11269__A2 (.I(_05524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11267__A2 (.I(_05524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11265__A2 (.I(_05524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11255__A2 (.I(_05524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11253__A2 (.I(_05524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11266__A2 (.I(_05527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11264__A2 (.I(_05527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11262__A2 (.I(_05527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11260__A2 (.I(_05527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11258__A2 (.I(_05527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11288__A2 (.I(_05534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11277__I (.I(_05534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11272__I (.I(_05534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11271__I (.I(_05534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11303__A2 (.I(_05547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11301__A2 (.I(_05547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11299__A2 (.I(_05547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11296__A2 (.I(_05547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11294__A2 (.I(_05547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11309__A2 (.I(_05548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11307__A2 (.I(_05548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11305__A2 (.I(_05548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11295__A2 (.I(_05548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11293__A2 (.I(_05548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11312__A2 (.I(_05558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11311__A2 (.I(_05558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(io_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(io_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout8_I (.I(\u_arbiter.i_wb_cpu_ack ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10573__A1 (.I(\u_arbiter.i_wb_cpu_ack ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10202__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10200__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05844__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10239__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10237__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05928__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10256__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10185__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05807__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10246__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10243__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05940__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10245__I (.I(\u_arbiter.i_wb_cpu_dbus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05945__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[22]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09605__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09600__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07012__I2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[30]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09628__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09624__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07012__I3 (.I(\u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[34]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09640__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09636__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[8]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09544__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09542__A3 (.I(\u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09533__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07705__A3 (.I(\u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[9]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09553__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09541__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07705__A4 (.I(\u_arbiter.i_wb_cpu_dbus_dat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[11]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09565__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09559__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07707__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06992__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[12]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09569__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07700__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[14]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09578__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09572__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07012__I1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07027__I (.I(\u_arbiter.i_wb_cpu_dbus_we ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06937__S (.I(\u_arbiter.i_wb_cpu_dbus_we ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06929__A1 (.I(\u_arbiter.i_wb_cpu_dbus_we ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06928__A1 (.I(\u_arbiter.i_wb_cpu_dbus_we ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06924__A1 (.I(\u_arbiter.i_wb_cpu_dbus_we ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07030__A1 (.I(\u_arbiter.i_wb_cpu_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07004__A1 (.I(\u_arbiter.i_wb_cpu_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05782__I (.I(\u_arbiter.i_wb_cpu_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10288__A1 (.I(\u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10286__B2 (.I(\u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09739__A2 (.I(\u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07695__A2 (.I(\u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05788__A1 (.I(\u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[3]_D  (.I(\u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10072__I1 (.I(\u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09712__I0 (.I(\u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09690__A2 (.I(\u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09531__A1 (.I(\u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[13]_D  (.I(\u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09893__I1 (.I(\u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09675__I0 (.I(\u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09585__A1 (.I(\u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[14]_D  (.I(\u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09984__I1 (.I(\u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09674__I0 (.I(\u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09588__A1 (.I(\u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[15]_D  (.I(\u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09989__A2 (.I(\u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09807__I0 (.I(\u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09686__A2 (.I(\u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09592__A1 (.I(\u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[16]_D  (.I(\u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10001__A2 (.I(\u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09752__I0 (.I(\u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09725__A2 (.I(\u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09596__A1 (.I(\u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[17]_D  (.I(\u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10011__I1 (.I(\u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09714__I0 (.I(\u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09706__A2 (.I(\u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09598__A1 (.I(\u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[18]_D  (.I(\u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10118__I1 (.I(\u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09716__A2 (.I(\u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09707__I0 (.I(\u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09601__A1 (.I(\u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[19]_D  (.I(\u_arbiter.i_wb_cpu_rdt[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10598__I0 (.I(\u_arbiter.i_wb_cpu_rdt[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10072__I0 (.I(\u_arbiter.i_wb_cpu_rdt[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09605__A1 (.I(\u_arbiter.i_wb_cpu_rdt[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[20]_D  (.I(\u_arbiter.i_wb_cpu_rdt[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10600__I0 (.I(\u_arbiter.i_wb_cpu_rdt[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10087__I0 (.I(\u_arbiter.i_wb_cpu_rdt[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09607__A1 (.I(\u_arbiter.i_wb_cpu_rdt[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[21]_D  (.I(\u_arbiter.i_wb_cpu_rdt[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10602__I0 (.I(\u_arbiter.i_wb_cpu_rdt[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10097__I0 (.I(\u_arbiter.i_wb_cpu_rdt[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09610__A1 (.I(\u_arbiter.i_wb_cpu_rdt[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[22]_D  (.I(\u_arbiter.i_wb_cpu_rdt[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10604__I0 (.I(\u_arbiter.i_wb_cpu_rdt[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10109__A2 (.I(\u_arbiter.i_wb_cpu_rdt[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09614__A1 (.I(\u_arbiter.i_wb_cpu_rdt[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[4]_D  (.I(\u_arbiter.i_wb_cpu_rdt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10087__I1 (.I(\u_arbiter.i_wb_cpu_rdt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09748__A2 (.I(\u_arbiter.i_wb_cpu_rdt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09693__I0 (.I(\u_arbiter.i_wb_cpu_rdt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09539__A1 (.I(\u_arbiter.i_wb_cpu_rdt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[23]_D  (.I(\u_arbiter.i_wb_cpu_rdt[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10606__I0 (.I(\u_arbiter.i_wb_cpu_rdt[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09826__I0 (.I(\u_arbiter.i_wb_cpu_rdt[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09617__A1 (.I(\u_arbiter.i_wb_cpu_rdt[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[24]_D  (.I(\u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10609__I0 (.I(\u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09843__I0 (.I(\u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09619__A1 (.I(\u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[25]_D  (.I(\u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10611__I0 (.I(\u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09859__I0 (.I(\u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09622__A1 (.I(\u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[26]_D  (.I(\u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10613__I0 (.I(\u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09936__I0 (.I(\u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09625__A1 (.I(\u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[27]_D  (.I(\u_arbiter.i_wb_cpu_rdt[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10615__I0 (.I(\u_arbiter.i_wb_cpu_rdt[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09952__I0 (.I(\u_arbiter.i_wb_cpu_rdt[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09627__A1 (.I(\u_arbiter.i_wb_cpu_rdt[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[28]_D  (.I(\u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10617__I0 (.I(\u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09968__A2 (.I(\u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09632__A1 (.I(\u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[29]_D  (.I(\u_arbiter.i_wb_cpu_rdt[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10620__I0 (.I(\u_arbiter.i_wb_cpu_rdt[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09893__I0 (.I(\u_arbiter.i_wb_cpu_rdt[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09634__A1 (.I(\u_arbiter.i_wb_cpu_rdt[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[30]_D  (.I(\u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10622__I0 (.I(\u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09984__I0 (.I(\u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09637__A1 (.I(\u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[31]_D  (.I(\u_arbiter.i_wb_cpu_rdt[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10624__I0 (.I(\u_arbiter.i_wb_cpu_rdt[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09990__A2 (.I(\u_arbiter.i_wb_cpu_rdt[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09640__A1 (.I(\u_arbiter.i_wb_cpu_rdt[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[32]_D  (.I(\u_arbiter.i_wb_cpu_rdt[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10626__I0 (.I(\u_arbiter.i_wb_cpu_rdt[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10002__A2 (.I(\u_arbiter.i_wb_cpu_rdt[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09643__A1 (.I(\u_arbiter.i_wb_cpu_rdt[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[5]_D  (.I(\u_arbiter.i_wb_cpu_rdt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10097__I1 (.I(\u_arbiter.i_wb_cpu_rdt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09702__I0 (.I(\u_arbiter.i_wb_cpu_rdt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09546__A1 (.I(\u_arbiter.i_wb_cpu_rdt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[33]_D  (.I(\u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10628__I0 (.I(\u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10011__I0 (.I(\u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09646__A1 (.I(\u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[34]_D  (.I(\u_arbiter.i_wb_cpu_rdt[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10630__I0 (.I(\u_arbiter.i_wb_cpu_rdt[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10118__I0 (.I(\u_arbiter.i_wb_cpu_rdt[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09648__A1 (.I(\u_arbiter.i_wb_cpu_rdt[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[7]_D  (.I(\u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09826__I1 (.I(\u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09701__I0 (.I(\u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09562__A1 (.I(\u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[8]_D  (.I(\u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09895__I0 (.I(\u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09843__I1 (.I(\u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09698__A2 (.I(\u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09564__A1 (.I(\u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[9]_D  (.I(\u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09859__I1 (.I(\u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09695__I0 (.I(\u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09569__A1 (.I(\u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[10]_D  (.I(\u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10027__A2 (.I(\u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09936__I1 (.I(\u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09677__I0 (.I(\u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09574__A1 (.I(\u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[11]_D  (.I(\u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09952__I1 (.I(\u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09729__I0 (.I(\u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09682__A2 (.I(\u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09578__A1 (.I(\u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[12]_D  (.I(\u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09995__A2 (.I(\u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09969__A2 (.I(\u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09676__I0 (.I(\u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09581__A1 (.I(\u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06981__A1 (.I(\u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06975__A1 (.I(\u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06974__A1 (.I(\u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06940__I (.I(\u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06925__A1 (.I(\u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06986__A1 (.I(\u_cpu.cpu.branch_op ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06930__A3 (.I(\u_cpu.cpu.branch_op ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06923__I (.I(\u_cpu.cpu.branch_op ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05728__A2 (.I(\u_cpu.cpu.branch_op ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05725__I (.I(\u_cpu.cpu.branch_op ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10571__A1 (.I(\u_cpu.cpu.bufreg.i_sh_signed ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10248__A1 (.I(\u_cpu.cpu.bufreg.i_sh_signed ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06924__A2 (.I(\u_cpu.cpu.bufreg.i_sh_signed ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09516__A1 (.I(\u_cpu.cpu.bufreg.lsb[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07012__S1 (.I(\u_cpu.cpu.bufreg.lsb[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05718__I (.I(\u_cpu.cpu.bufreg.lsb[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06961__I (.I(\u_cpu.cpu.bufreg2.i_cnt_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06932__A1 (.I(\u_cpu.cpu.bufreg2.i_cnt_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06931__A1 (.I(\u_cpu.cpu.bufreg2.i_cnt_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10056__A1 (.I(\u_cpu.cpu.csr_imm ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05740__I (.I(\u_cpu.cpu.csr_imm ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11120__A1 (.I(\u_cpu.cpu.ctrl.i_iscomp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07002__A2 (.I(\u_cpu.cpu.ctrl.i_iscomp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07001__A2 (.I(\u_cpu.cpu.ctrl.i_iscomp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10346__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10343__B2 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05926__A2 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05921__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05918__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10356__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10354__B2 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05942__I (.I(\u_cpu.cpu.ctrl.o_ibus_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05939__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10300__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10298__B2 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05834__A2 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05825__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05824__B (.I(\u_cpu.cpu.ctrl.o_ibus_adr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10302__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10300__B2 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05834__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05829__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11111__A1 (.I(\u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06964__A2 (.I(\u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05763__A2 (.I(\u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05731__I (.I(\u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06963__I (.I(\u_cpu.cpu.decode.op21 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05744__A1 (.I(\u_cpu.cpu.decode.op21 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05733__A3 (.I(\u_cpu.cpu.decode.op21 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05732__A1 (.I(\u_cpu.cpu.decode.op21 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05727__A1 (.I(\u_cpu.cpu.decode.op21 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07028__A2 (.I(\u_cpu.cpu.decode.opcode[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07007__I (.I(\u_cpu.cpu.decode.opcode[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06986__A2 (.I(\u_cpu.cpu.decode.opcode[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06927__A3 (.I(\u_cpu.cpu.decode.opcode[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06930__A2 (.I(\u_cpu.cpu.decode.opcode[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06927__A1 (.I(\u_cpu.cpu.decode.opcode[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05728__A1 (.I(\u_cpu.cpu.decode.opcode[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05723__I (.I(\u_cpu.cpu.decode.opcode[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05820__A1 (.I(\u_cpu.cpu.genblk1.align.ctrl_misal ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05790__I (.I(\u_cpu.cpu.genblk1.align.ctrl_misal ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10624__I1 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09807__I1 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09685__A2 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10609__I1 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09895__I1 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09697__A2 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10611__I1 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09695__I1 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10613__I1 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10026__A2 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09677__I1 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10617__I1 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09994__A2 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09676__I1 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[1]_D  (.I(\u_cpu.cpu.genblk3.csr.i_mtip ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10123__A3 (.I(\u_cpu.cpu.genblk3.csr.i_mtip ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11118__A1 (.I(\u_cpu.cpu.genblk3.csr.mstatus_mie ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11108__I0 (.I(\u_cpu.cpu.genblk3.csr.mstatus_mie ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10123__A2 (.I(\u_cpu.cpu.genblk3.csr.mstatus_mie ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06967__B2 (.I(\u_cpu.cpu.genblk3.csr.mstatus_mie ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10455__I0 (.I(\u_cpu.cpu.immdec.imm11_7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10446__A1 (.I(\u_cpu.cpu.immdec.imm11_7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07131__A1 (.I(\u_cpu.cpu.immdec.imm11_7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07116__A1 (.I(\u_cpu.cpu.immdec.imm11_7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07213__I (.I(\u_cpu.cpu.immdec.imm11_7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07147__A1 (.I(\u_cpu.cpu.immdec.imm11_7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07120__A1 (.I(\u_cpu.cpu.immdec.imm11_7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10112__A2 (.I(\u_cpu.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09927__A1 (.I(\u_cpu.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06929__B (.I(\u_cpu.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05739__A1 (.I(\u_cpu.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09932__I (.I(\u_cpu.cpu.immdec.imm24_20[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09930__B2 (.I(\u_cpu.cpu.immdec.imm24_20[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05774__A1 (.I(\u_cpu.cpu.immdec.imm24_20[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09956__A1 (.I(\u_cpu.cpu.immdec.imm24_20[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09946__A1 (.I(\u_cpu.cpu.immdec.imm24_20[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05752__A1 (.I(\u_cpu.cpu.immdec.imm24_20[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09976__A1 (.I(\u_cpu.cpu.immdec.imm30_25[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09971__A1 (.I(\u_cpu.cpu.immdec.imm30_25[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10119__A1 (.I(\u_cpu.cpu.immdec.imm31 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07019__A1 (.I(\u_cpu.cpu.immdec.imm31 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06931__A2 (.I(\u_cpu.cpu.immdec.imm31 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09128__I (.I(\u_cpu.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07022__A2 (.I(\u_cpu.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07011__B1 (.I(\u_cpu.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06956__A3 (.I(\u_cpu.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12690__D (.I(\u_cpu.cpu.o_wdata0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07337__I1 (.I(\u_cpu.cpu.o_wdata0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07201__A2 (.I(\u_cpu.cpu.o_wdata0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12704__D (.I(\u_cpu.cpu.o_wdata1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09196__A1 (.I(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07697__A1 (.I(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05743__A2 (.I(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05735__I (.I(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10252__A2 (.I(\u_cpu.cpu.state.o_cnt_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07082__A2 (.I(\u_cpu.cpu.state.o_cnt_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07000__I (.I(\u_cpu.cpu.state.o_cnt_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06918__A2 (.I(\u_cpu.cpu.state.o_cnt_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07207__A1 (.I(\u_cpu.raddr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06041__I (.I(\u_cpu.raddr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06006__I (.I(\u_cpu.raddr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05958__I (.I(\u_cpu.raddr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11258__A1 (.I(\u_cpu.rf_ram.memory[100][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06394__I0 (.I(\u_cpu.rf_ram.memory[100][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10663__A1 (.I(\u_cpu.rf_ram.memory[102][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06109__I2 (.I(\u_cpu.rf_ram.memory[102][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10665__A1 (.I(\u_cpu.rf_ram.memory[102][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06280__I2 (.I(\u_cpu.rf_ram.memory[102][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10668__A1 (.I(\u_cpu.rf_ram.memory[102][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06394__I2 (.I(\u_cpu.rf_ram.memory[102][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10670__A1 (.I(\u_cpu.rf_ram.memory[102][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06509__I2 (.I(\u_cpu.rf_ram.memory[102][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10672__A1 (.I(\u_cpu.rf_ram.memory[102][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06608__I2 (.I(\u_cpu.rf_ram.memory[102][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10704__A1 (.I(\u_cpu.rf_ram.memory[104][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06105__I0 (.I(\u_cpu.rf_ram.memory[104][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10706__A1 (.I(\u_cpu.rf_ram.memory[104][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06277__I0 (.I(\u_cpu.rf_ram.memory[104][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10717__A1 (.I(\u_cpu.rf_ram.memory[104][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06782__I0 (.I(\u_cpu.rf_ram.memory[104][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10719__A1 (.I(\u_cpu.rf_ram.memory[104][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06870__I0 (.I(\u_cpu.rf_ram.memory[104][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10801__A1 (.I(\u_cpu.rf_ram.memory[106][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06606__I2 (.I(\u_cpu.rf_ram.memory[106][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10864__A1 (.I(\u_cpu.rf_ram.memory[108][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06504__I0 (.I(\u_cpu.rf_ram.memory[108][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10867__A1 (.I(\u_cpu.rf_ram.memory[108][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06604__I0 (.I(\u_cpu.rf_ram.memory[108][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10870__A1 (.I(\u_cpu.rf_ram.memory[108][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06692__I0 (.I(\u_cpu.rf_ram.memory[108][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10370__A1 (.I(\u_cpu.rf_ram.memory[109][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06101__I1 (.I(\u_cpu.rf_ram.memory[109][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10372__A1 (.I(\u_cpu.rf_ram.memory[109][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06274__I1 (.I(\u_cpu.rf_ram.memory[109][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10381__A1 (.I(\u_cpu.rf_ram.memory[109][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06692__I1 (.I(\u_cpu.rf_ram.memory[109][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10385__A1 (.I(\u_cpu.rf_ram.memory[109][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06868__I1 (.I(\u_cpu.rf_ram.memory[109][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10981__A1 (.I(\u_cpu.rf_ram.memory[110][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06101__I2 (.I(\u_cpu.rf_ram.memory[110][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10988__A1 (.I(\u_cpu.rf_ram.memory[110][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06387__I2 (.I(\u_cpu.rf_ram.memory[110][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09415__A1 (.I(\u_cpu.rf_ram.memory[112][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06405__I0 (.I(\u_cpu.rf_ram.memory[112][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09417__A1 (.I(\u_cpu.rf_ram.memory[112][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06520__I0 (.I(\u_cpu.rf_ram.memory[112][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09419__A1 (.I(\u_cpu.rf_ram.memory[112][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06617__I0 (.I(\u_cpu.rf_ram.memory[112][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09421__A1 (.I(\u_cpu.rf_ram.memory[112][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06705__I0 (.I(\u_cpu.rf_ram.memory[112][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09423__A1 (.I(\u_cpu.rf_ram.memory[112][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06793__I0 (.I(\u_cpu.rf_ram.memory[112][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09425__A1 (.I(\u_cpu.rf_ram.memory[112][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06881__I0 (.I(\u_cpu.rf_ram.memory[112][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09876__A1 (.I(\u_cpu.rf_ram.memory[114][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06132__I2 (.I(\u_cpu.rf_ram.memory[114][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09878__A1 (.I(\u_cpu.rf_ram.memory[114][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06293__I2 (.I(\u_cpu.rf_ram.memory[114][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09881__A1 (.I(\u_cpu.rf_ram.memory[114][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06405__I2 (.I(\u_cpu.rf_ram.memory[114][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09883__A1 (.I(\u_cpu.rf_ram.memory[114][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06520__I2 (.I(\u_cpu.rf_ram.memory[114][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09889__A1 (.I(\u_cpu.rf_ram.memory[114][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06793__I2 (.I(\u_cpu.rf_ram.memory[114][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09891__A1 (.I(\u_cpu.rf_ram.memory[114][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06881__I2 (.I(\u_cpu.rf_ram.memory[114][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09479__A1 (.I(\u_cpu.rf_ram.memory[116][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06137__I0 (.I(\u_cpu.rf_ram.memory[116][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09481__A1 (.I(\u_cpu.rf_ram.memory[116][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06295__I0 (.I(\u_cpu.rf_ram.memory[116][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09278__A1 (.I(\u_cpu.rf_ram.memory[117][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06137__I1 (.I(\u_cpu.rf_ram.memory[117][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09280__A1 (.I(\u_cpu.rf_ram.memory[117][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06295__I1 (.I(\u_cpu.rf_ram.memory[117][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09287__A1 (.I(\u_cpu.rf_ram.memory[117][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06619__I1 (.I(\u_cpu.rf_ram.memory[117][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09289__A1 (.I(\u_cpu.rf_ram.memory[117][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06707__I1 (.I(\u_cpu.rf_ram.memory[117][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09291__A1 (.I(\u_cpu.rf_ram.memory[117][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06795__I1 (.I(\u_cpu.rf_ram.memory[117][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09293__A1 (.I(\u_cpu.rf_ram.memory[117][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06883__I1 (.I(\u_cpu.rf_ram.memory[117][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09326__A1 (.I(\u_cpu.rf_ram.memory[118][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06137__I2 (.I(\u_cpu.rf_ram.memory[118][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09328__A1 (.I(\u_cpu.rf_ram.memory[118][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06295__I2 (.I(\u_cpu.rf_ram.memory[118][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09331__A1 (.I(\u_cpu.rf_ram.memory[118][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06407__I2 (.I(\u_cpu.rf_ram.memory[118][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09333__A1 (.I(\u_cpu.rf_ram.memory[118][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06523__I2 (.I(\u_cpu.rf_ram.memory[118][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09335__A1 (.I(\u_cpu.rf_ram.memory[118][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06619__I2 (.I(\u_cpu.rf_ram.memory[118][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09337__A1 (.I(\u_cpu.rf_ram.memory[118][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06707__I2 (.I(\u_cpu.rf_ram.memory[118][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09339__A1 (.I(\u_cpu.rf_ram.memory[118][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06795__I2 (.I(\u_cpu.rf_ram.memory[118][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09341__A1 (.I(\u_cpu.rf_ram.memory[118][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06883__I2 (.I(\u_cpu.rf_ram.memory[118][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07792__A1 (.I(\u_cpu.rf_ram.memory[119][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06137__I3 (.I(\u_cpu.rf_ram.memory[119][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07795__A1 (.I(\u_cpu.rf_ram.memory[119][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06295__I3 (.I(\u_cpu.rf_ram.memory[119][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07799__A1 (.I(\u_cpu.rf_ram.memory[119][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06407__I3 (.I(\u_cpu.rf_ram.memory[119][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07802__A1 (.I(\u_cpu.rf_ram.memory[119][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06523__I3 (.I(\u_cpu.rf_ram.memory[119][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07805__A1 (.I(\u_cpu.rf_ram.memory[119][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06619__I3 (.I(\u_cpu.rf_ram.memory[119][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07808__A1 (.I(\u_cpu.rf_ram.memory[119][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06707__I3 (.I(\u_cpu.rf_ram.memory[119][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07811__A1 (.I(\u_cpu.rf_ram.memory[119][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06795__I3 (.I(\u_cpu.rf_ram.memory[119][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07814__A1 (.I(\u_cpu.rf_ram.memory[119][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06883__I3 (.I(\u_cpu.rf_ram.memory[119][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09315__A1 (.I(\u_cpu.rf_ram.memory[120][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06703__I0 (.I(\u_cpu.rf_ram.memory[120][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09357__A1 (.I(\u_cpu.rf_ram.memory[121][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06703__I1 (.I(\u_cpu.rf_ram.memory[121][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09040__A1 (.I(\u_cpu.rf_ram.memory[123][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06290__I3 (.I(\u_cpu.rf_ram.memory[123][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09044__A1 (.I(\u_cpu.rf_ram.memory[123][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06403__I3 (.I(\u_cpu.rf_ram.memory[123][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09047__A1 (.I(\u_cpu.rf_ram.memory[123][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06517__I3 (.I(\u_cpu.rf_ram.memory[123][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09050__A1 (.I(\u_cpu.rf_ram.memory[123][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06615__I3 (.I(\u_cpu.rf_ram.memory[123][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09024__A1 (.I(\u_cpu.rf_ram.memory[124][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06613__I0 (.I(\u_cpu.rf_ram.memory[124][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08995__A1 (.I(\u_cpu.rf_ram.memory[125][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06121__I1 (.I(\u_cpu.rf_ram.memory[125][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08997__A1 (.I(\u_cpu.rf_ram.memory[125][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06286__I1 (.I(\u_cpu.rf_ram.memory[125][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09000__A1 (.I(\u_cpu.rf_ram.memory[125][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06401__I1 (.I(\u_cpu.rf_ram.memory[125][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09002__A1 (.I(\u_cpu.rf_ram.memory[125][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06515__I1 (.I(\u_cpu.rf_ram.memory[125][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09004__A1 (.I(\u_cpu.rf_ram.memory[125][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06613__I1 (.I(\u_cpu.rf_ram.memory[125][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09008__A1 (.I(\u_cpu.rf_ram.memory[125][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06789__I1 (.I(\u_cpu.rf_ram.memory[125][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08921__A1 (.I(\u_cpu.rf_ram.memory[128][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06211__I0 (.I(\u_cpu.rf_ram.memory[128][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08930__A1 (.I(\u_cpu.rf_ram.memory[128][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06443__I0 (.I(\u_cpu.rf_ram.memory[128][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08934__A1 (.I(\u_cpu.rf_ram.memory[128][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06558__I0 (.I(\u_cpu.rf_ram.memory[128][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07821__A1 (.I(\u_cpu.rf_ram.memory[129][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06211__I1 (.I(\u_cpu.rf_ram.memory[129][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07823__A1 (.I(\u_cpu.rf_ram.memory[129][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06332__I1 (.I(\u_cpu.rf_ram.memory[129][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07826__A1 (.I(\u_cpu.rf_ram.memory[129][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06443__I1 (.I(\u_cpu.rf_ram.memory[129][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07828__A1 (.I(\u_cpu.rf_ram.memory[129][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06558__I1 (.I(\u_cpu.rf_ram.memory[129][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07830__A1 (.I(\u_cpu.rf_ram.memory[129][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06647__I1 (.I(\u_cpu.rf_ram.memory[129][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07832__A1 (.I(\u_cpu.rf_ram.memory[129][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06735__I1 (.I(\u_cpu.rf_ram.memory[129][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07834__A1 (.I(\u_cpu.rf_ram.memory[129][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06823__I1 (.I(\u_cpu.rf_ram.memory[129][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07836__A1 (.I(\u_cpu.rf_ram.memory[129][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06911__I1 (.I(\u_cpu.rf_ram.memory[129][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08731__A1 (.I(\u_cpu.rf_ram.memory[136][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06200__I0 (.I(\u_cpu.rf_ram.memory[136][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08733__A1 (.I(\u_cpu.rf_ram.memory[136][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06327__I0 (.I(\u_cpu.rf_ram.memory[136][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08736__A1 (.I(\u_cpu.rf_ram.memory[136][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06439__I0 (.I(\u_cpu.rf_ram.memory[136][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08738__A1 (.I(\u_cpu.rf_ram.memory[136][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06553__I0 (.I(\u_cpu.rf_ram.memory[136][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08740__A1 (.I(\u_cpu.rf_ram.memory[136][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06643__I0 (.I(\u_cpu.rf_ram.memory[136][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08742__A1 (.I(\u_cpu.rf_ram.memory[136][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06731__I0 (.I(\u_cpu.rf_ram.memory[136][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08744__A1 (.I(\u_cpu.rf_ram.memory[136][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06819__I0 (.I(\u_cpu.rf_ram.memory[136][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08746__A1 (.I(\u_cpu.rf_ram.memory[136][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06907__I0 (.I(\u_cpu.rf_ram.memory[136][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08691__A1 (.I(\u_cpu.rf_ram.memory[137][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06439__I1 (.I(\u_cpu.rf_ram.memory[137][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08694__A1 (.I(\u_cpu.rf_ram.memory[137][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06553__I1 (.I(\u_cpu.rf_ram.memory[137][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08700__A1 (.I(\u_cpu.rf_ram.memory[137][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06731__I1 (.I(\u_cpu.rf_ram.memory[137][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08703__A1 (.I(\u_cpu.rf_ram.memory[137][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06819__I1 (.I(\u_cpu.rf_ram.memory[137][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08706__A1 (.I(\u_cpu.rf_ram.memory[137][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06907__I1 (.I(\u_cpu.rf_ram.memory[137][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08643__A1 (.I(\u_cpu.rf_ram.memory[138][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06200__I2 (.I(\u_cpu.rf_ram.memory[138][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08645__A1 (.I(\u_cpu.rf_ram.memory[138][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06327__I2 (.I(\u_cpu.rf_ram.memory[138][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08648__A1 (.I(\u_cpu.rf_ram.memory[138][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06439__I2 (.I(\u_cpu.rf_ram.memory[138][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08650__A1 (.I(\u_cpu.rf_ram.memory[138][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06553__I2 (.I(\u_cpu.rf_ram.memory[138][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08652__A1 (.I(\u_cpu.rf_ram.memory[138][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06643__I2 (.I(\u_cpu.rf_ram.memory[138][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08658__A1 (.I(\u_cpu.rf_ram.memory[138][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06907__I2 (.I(\u_cpu.rf_ram.memory[138][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08616__A1 (.I(\u_cpu.rf_ram.memory[143][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06733__I3 (.I(\u_cpu.rf_ram.memory[143][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08618__A1 (.I(\u_cpu.rf_ram.memory[143][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06821__I3 (.I(\u_cpu.rf_ram.memory[143][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08620__A1 (.I(\u_cpu.rf_ram.memory[143][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06909__I3 (.I(\u_cpu.rf_ram.memory[143][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07754__A1 (.I(\u_cpu.rf_ram.memory[17][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06468__I1 (.I(\u_cpu.rf_ram.memory[17][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07264__A1 (.I(\u_cpu.rf_ram.memory[18][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06237__I2 (.I(\u_cpu.rf_ram.memory[18][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07267__A1 (.I(\u_cpu.rf_ram.memory[18][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06354__I2 (.I(\u_cpu.rf_ram.memory[18][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07269__A1 (.I(\u_cpu.rf_ram.memory[18][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06468__I2 (.I(\u_cpu.rf_ram.memory[18][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07271__A1 (.I(\u_cpu.rf_ram.memory[18][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06577__I2 (.I(\u_cpu.rf_ram.memory[18][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07273__A1 (.I(\u_cpu.rf_ram.memory[18][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06665__I2 (.I(\u_cpu.rf_ram.memory[18][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07275__A1 (.I(\u_cpu.rf_ram.memory[18][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06753__I2 (.I(\u_cpu.rf_ram.memory[18][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08192__A1 (.I(\u_cpu.rf_ram.memory[19][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06009__I3 (.I(\u_cpu.rf_ram.memory[19][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08194__A1 (.I(\u_cpu.rf_ram.memory[19][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06237__I3 (.I(\u_cpu.rf_ram.memory[19][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08197__A1 (.I(\u_cpu.rf_ram.memory[19][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06354__I3 (.I(\u_cpu.rf_ram.memory[19][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08199__A1 (.I(\u_cpu.rf_ram.memory[19][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06468__I3 (.I(\u_cpu.rf_ram.memory[19][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08201__A1 (.I(\u_cpu.rf_ram.memory[19][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06577__I3 (.I(\u_cpu.rf_ram.memory[19][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08203__A1 (.I(\u_cpu.rf_ram.memory[19][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06665__I3 (.I(\u_cpu.rf_ram.memory[19][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08205__A1 (.I(\u_cpu.rf_ram.memory[19][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06753__I3 (.I(\u_cpu.rf_ram.memory[19][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08207__A1 (.I(\u_cpu.rf_ram.memory[19][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06841__I3 (.I(\u_cpu.rf_ram.memory[19][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07285__A1 (.I(\u_cpu.rf_ram.memory[20][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06000__I0 (.I(\u_cpu.rf_ram.memory[20][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07287__A1 (.I(\u_cpu.rf_ram.memory[20][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06234__I0 (.I(\u_cpu.rf_ram.memory[20][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07290__A1 (.I(\u_cpu.rf_ram.memory[20][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06351__I0 (.I(\u_cpu.rf_ram.memory[20][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07292__A1 (.I(\u_cpu.rf_ram.memory[20][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06465__I0 (.I(\u_cpu.rf_ram.memory[20][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07294__A1 (.I(\u_cpu.rf_ram.memory[20][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06575__I0 (.I(\u_cpu.rf_ram.memory[20][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07296__A1 (.I(\u_cpu.rf_ram.memory[20][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06663__I0 (.I(\u_cpu.rf_ram.memory[20][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07298__A1 (.I(\u_cpu.rf_ram.memory[20][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06751__I0 (.I(\u_cpu.rf_ram.memory[20][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07300__A1 (.I(\u_cpu.rf_ram.memory[20][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06839__I0 (.I(\u_cpu.rf_ram.memory[20][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07220__A1 (.I(\u_cpu.rf_ram.memory[21][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06000__I1 (.I(\u_cpu.rf_ram.memory[21][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07222__A1 (.I(\u_cpu.rf_ram.memory[21][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06234__I1 (.I(\u_cpu.rf_ram.memory[21][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07225__A1 (.I(\u_cpu.rf_ram.memory[21][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06351__I1 (.I(\u_cpu.rf_ram.memory[21][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07227__A1 (.I(\u_cpu.rf_ram.memory[21][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06465__I1 (.I(\u_cpu.rf_ram.memory[21][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07229__A1 (.I(\u_cpu.rf_ram.memory[21][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06575__I1 (.I(\u_cpu.rf_ram.memory[21][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07235__A1 (.I(\u_cpu.rf_ram.memory[21][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06839__I1 (.I(\u_cpu.rf_ram.memory[21][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08899__A1 (.I(\u_cpu.rf_ram.memory[22][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06000__I2 (.I(\u_cpu.rf_ram.memory[22][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08901__A1 (.I(\u_cpu.rf_ram.memory[22][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06234__I2 (.I(\u_cpu.rf_ram.memory[22][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08904__A1 (.I(\u_cpu.rf_ram.memory[22][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06351__I2 (.I(\u_cpu.rf_ram.memory[22][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08906__A1 (.I(\u_cpu.rf_ram.memory[22][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06465__I2 (.I(\u_cpu.rf_ram.memory[22][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08908__A1 (.I(\u_cpu.rf_ram.memory[22][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06575__I2 (.I(\u_cpu.rf_ram.memory[22][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08910__A1 (.I(\u_cpu.rf_ram.memory[22][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06663__I2 (.I(\u_cpu.rf_ram.memory[22][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08912__A1 (.I(\u_cpu.rf_ram.memory[22][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06751__I2 (.I(\u_cpu.rf_ram.memory[22][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08914__A1 (.I(\u_cpu.rf_ram.memory[22][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06839__I2 (.I(\u_cpu.rf_ram.memory[22][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11300__A1 (.I(\u_cpu.rf_ram.memory[23][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06465__I3 (.I(\u_cpu.rf_ram.memory[23][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11302__A1 (.I(\u_cpu.rf_ram.memory[23][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06575__I3 (.I(\u_cpu.rf_ram.memory[23][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11155__A1 (.I(\u_cpu.rf_ram.memory[26][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06026__I2 (.I(\u_cpu.rf_ram.memory[26][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11128__A1 (.I(\u_cpu.rf_ram.memory[27][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06026__I3 (.I(\u_cpu.rf_ram.memory[27][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11131__A1 (.I(\u_cpu.rf_ram.memory[27][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06242__I3 (.I(\u_cpu.rf_ram.memory[27][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11138__A1 (.I(\u_cpu.rf_ram.memory[27][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06473__I3 (.I(\u_cpu.rf_ram.memory[27][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11141__A1 (.I(\u_cpu.rf_ram.memory[27][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06581__I3 (.I(\u_cpu.rf_ram.memory[27][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11144__A1 (.I(\u_cpu.rf_ram.memory[27][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06669__I3 (.I(\u_cpu.rf_ram.memory[27][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11147__A1 (.I(\u_cpu.rf_ram.memory[27][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06757__I3 (.I(\u_cpu.rf_ram.memory[27][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11150__A1 (.I(\u_cpu.rf_ram.memory[27][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06845__I3 (.I(\u_cpu.rf_ram.memory[27][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10580__A1 (.I(\u_cpu.rf_ram.memory[28][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06018__I0 (.I(\u_cpu.rf_ram.memory[28][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10582__A1 (.I(\u_cpu.rf_ram.memory[28][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06239__I0 (.I(\u_cpu.rf_ram.memory[28][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10585__A1 (.I(\u_cpu.rf_ram.memory[28][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06357__I0 (.I(\u_cpu.rf_ram.memory[28][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10587__A1 (.I(\u_cpu.rf_ram.memory[28][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06471__I0 (.I(\u_cpu.rf_ram.memory[28][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10589__A1 (.I(\u_cpu.rf_ram.memory[28][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06579__I0 (.I(\u_cpu.rf_ram.memory[28][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10593__A1 (.I(\u_cpu.rf_ram.memory[28][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06755__I0 (.I(\u_cpu.rf_ram.memory[28][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10595__A1 (.I(\u_cpu.rf_ram.memory[28][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06843__I0 (.I(\u_cpu.rf_ram.memory[28][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08082__A1 (.I(\u_cpu.rf_ram.memory[29][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06018__I1 (.I(\u_cpu.rf_ram.memory[29][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08084__A1 (.I(\u_cpu.rf_ram.memory[29][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06239__I1 (.I(\u_cpu.rf_ram.memory[29][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08091__A1 (.I(\u_cpu.rf_ram.memory[29][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06579__I1 (.I(\u_cpu.rf_ram.memory[29][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08093__A1 (.I(\u_cpu.rf_ram.memory[29][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06667__I1 (.I(\u_cpu.rf_ram.memory[29][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08095__A1 (.I(\u_cpu.rf_ram.memory[29][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06755__I1 (.I(\u_cpu.rf_ram.memory[29][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08097__A1 (.I(\u_cpu.rf_ram.memory[29][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06843__I1 (.I(\u_cpu.rf_ram.memory[29][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10130__A1 (.I(\u_cpu.rf_ram.memory[32][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06091__I0 (.I(\u_cpu.rf_ram.memory[32][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10134__A1 (.I(\u_cpu.rf_ram.memory[32][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06269__I0 (.I(\u_cpu.rf_ram.memory[32][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10139__A1 (.I(\u_cpu.rf_ram.memory[32][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06380__I0 (.I(\u_cpu.rf_ram.memory[32][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10143__A1 (.I(\u_cpu.rf_ram.memory[32][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06498__I0 (.I(\u_cpu.rf_ram.memory[32][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10147__A1 (.I(\u_cpu.rf_ram.memory[32][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06599__I0 (.I(\u_cpu.rf_ram.memory[32][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10151__A1 (.I(\u_cpu.rf_ram.memory[32][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06687__I0 (.I(\u_cpu.rf_ram.memory[32][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10155__A1 (.I(\u_cpu.rf_ram.memory[32][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06775__I0 (.I(\u_cpu.rf_ram.memory[32][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10159__A1 (.I(\u_cpu.rf_ram.memory[32][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06863__I0 (.I(\u_cpu.rf_ram.memory[32][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09504__A1 (.I(\u_cpu.rf_ram.memory[33][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06380__I1 (.I(\u_cpu.rf_ram.memory[33][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09506__A1 (.I(\u_cpu.rf_ram.memory[33][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06498__I1 (.I(\u_cpu.rf_ram.memory[33][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09508__A1 (.I(\u_cpu.rf_ram.memory[33][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06599__I1 (.I(\u_cpu.rf_ram.memory[33][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09510__A1 (.I(\u_cpu.rf_ram.memory[33][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06687__I1 (.I(\u_cpu.rf_ram.memory[33][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09512__A1 (.I(\u_cpu.rf_ram.memory[33][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06775__I1 (.I(\u_cpu.rf_ram.memory[33][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09514__A1 (.I(\u_cpu.rf_ram.memory[33][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06863__I1 (.I(\u_cpu.rf_ram.memory[33][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09260__A1 (.I(\u_cpu.rf_ram.memory[34][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06269__I2 (.I(\u_cpu.rf_ram.memory[34][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09104__A1 (.I(\u_cpu.rf_ram.memory[36][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06083__I0 (.I(\u_cpu.rf_ram.memory[36][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09106__A1 (.I(\u_cpu.rf_ram.memory[36][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06267__I0 (.I(\u_cpu.rf_ram.memory[36][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09109__A1 (.I(\u_cpu.rf_ram.memory[36][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06376__I0 (.I(\u_cpu.rf_ram.memory[36][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09111__A1 (.I(\u_cpu.rf_ram.memory[36][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06496__I0 (.I(\u_cpu.rf_ram.memory[36][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09113__A1 (.I(\u_cpu.rf_ram.memory[36][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06597__I0 (.I(\u_cpu.rf_ram.memory[36][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09115__A1 (.I(\u_cpu.rf_ram.memory[36][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06685__I0 (.I(\u_cpu.rf_ram.memory[36][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09117__A1 (.I(\u_cpu.rf_ram.memory[36][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06773__I0 (.I(\u_cpu.rf_ram.memory[36][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09119__A1 (.I(\u_cpu.rf_ram.memory[36][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06861__I0 (.I(\u_cpu.rf_ram.memory[36][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09086__A1 (.I(\u_cpu.rf_ram.memory[37][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06267__I1 (.I(\u_cpu.rf_ram.memory[37][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09089__A1 (.I(\u_cpu.rf_ram.memory[37][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06376__I1 (.I(\u_cpu.rf_ram.memory[37][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09097__A1 (.I(\u_cpu.rf_ram.memory[37][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06773__I1 (.I(\u_cpu.rf_ram.memory[37][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08663__A1 (.I(\u_cpu.rf_ram.memory[39][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06083__I3 (.I(\u_cpu.rf_ram.memory[39][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08665__A1 (.I(\u_cpu.rf_ram.memory[39][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06267__I3 (.I(\u_cpu.rf_ram.memory[39][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08668__A1 (.I(\u_cpu.rf_ram.memory[39][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06376__I3 (.I(\u_cpu.rf_ram.memory[39][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08670__A1 (.I(\u_cpu.rf_ram.memory[39][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06496__I3 (.I(\u_cpu.rf_ram.memory[39][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08672__A1 (.I(\u_cpu.rf_ram.memory[39][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06597__I3 (.I(\u_cpu.rf_ram.memory[39][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08674__A1 (.I(\u_cpu.rf_ram.memory[39][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06685__I3 (.I(\u_cpu.rf_ram.memory[39][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08676__A1 (.I(\u_cpu.rf_ram.memory[39][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06773__I3 (.I(\u_cpu.rf_ram.memory[39][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08678__A1 (.I(\u_cpu.rf_ram.memory[39][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06861__I3 (.I(\u_cpu.rf_ram.memory[39][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07771__A1 (.I(\u_cpu.rf_ram.memory[40][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06261__I0 (.I(\u_cpu.rf_ram.memory[40][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07776__A1 (.I(\u_cpu.rf_ram.memory[40][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06490__I0 (.I(\u_cpu.rf_ram.memory[40][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07780__A1 (.I(\u_cpu.rf_ram.memory[40][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06681__I0 (.I(\u_cpu.rf_ram.memory[40][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07782__A1 (.I(\u_cpu.rf_ram.memory[40][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06769__I0 (.I(\u_cpu.rf_ram.memory[40][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07554__A1 (.I(\u_cpu.rf_ram.memory[41][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06072__I1 (.I(\u_cpu.rf_ram.memory[41][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07556__A1 (.I(\u_cpu.rf_ram.memory[41][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06261__I1 (.I(\u_cpu.rf_ram.memory[41][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07559__A1 (.I(\u_cpu.rf_ram.memory[41][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06371__I1 (.I(\u_cpu.rf_ram.memory[41][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07561__A1 (.I(\u_cpu.rf_ram.memory[41][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06490__I1 (.I(\u_cpu.rf_ram.memory[41][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07563__A1 (.I(\u_cpu.rf_ram.memory[41][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06593__I1 (.I(\u_cpu.rf_ram.memory[41][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07565__A1 (.I(\u_cpu.rf_ram.memory[41][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06681__I1 (.I(\u_cpu.rf_ram.memory[41][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07567__A1 (.I(\u_cpu.rf_ram.memory[41][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06769__I1 (.I(\u_cpu.rf_ram.memory[41][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07569__A1 (.I(\u_cpu.rf_ram.memory[41][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06857__I1 (.I(\u_cpu.rf_ram.memory[41][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07445__A1 (.I(\u_cpu.rf_ram.memory[42][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06681__I2 (.I(\u_cpu.rf_ram.memory[42][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07500__A1 (.I(\u_cpu.rf_ram.memory[44][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06077__I0 (.I(\u_cpu.rf_ram.memory[44][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07503__A1 (.I(\u_cpu.rf_ram.memory[44][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06264__I0 (.I(\u_cpu.rf_ram.memory[44][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07459__A1 (.I(\u_cpu.rf_ram.memory[46][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06374__I2 (.I(\u_cpu.rf_ram.memory[46][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07463__A1 (.I(\u_cpu.rf_ram.memory[46][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06595__I2 (.I(\u_cpu.rf_ram.memory[46][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07465__A1 (.I(\u_cpu.rf_ram.memory[46][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06683__I2 (.I(\u_cpu.rf_ram.memory[46][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07620__A1 (.I(\u_cpu.rf_ram.memory[47][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06077__I3 (.I(\u_cpu.rf_ram.memory[47][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07624__A1 (.I(\u_cpu.rf_ram.memory[47][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06264__I3 (.I(\u_cpu.rf_ram.memory[47][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07637__A1 (.I(\u_cpu.rf_ram.memory[47][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06595__I3 (.I(\u_cpu.rf_ram.memory[47][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07641__A1 (.I(\u_cpu.rf_ram.memory[47][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06683__I3 (.I(\u_cpu.rf_ram.memory[47][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07645__A1 (.I(\u_cpu.rf_ram.memory[47][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06771__I3 (.I(\u_cpu.rf_ram.memory[47][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07649__A1 (.I(\u_cpu.rf_ram.memory[47][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06859__I3 (.I(\u_cpu.rf_ram.memory[47][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08711__A1 (.I(\u_cpu.rf_ram.memory[49][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06044__I1 (.I(\u_cpu.rf_ram.memory[49][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08713__A1 (.I(\u_cpu.rf_ram.memory[49][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06250__I1 (.I(\u_cpu.rf_ram.memory[49][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08716__A1 (.I(\u_cpu.rf_ram.memory[49][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06364__I1 (.I(\u_cpu.rf_ram.memory[49][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08718__A1 (.I(\u_cpu.rf_ram.memory[49][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06479__I1 (.I(\u_cpu.rf_ram.memory[49][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08720__A1 (.I(\u_cpu.rf_ram.memory[49][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06586__I1 (.I(\u_cpu.rf_ram.memory[49][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08722__A1 (.I(\u_cpu.rf_ram.memory[49][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06674__I1 (.I(\u_cpu.rf_ram.memory[49][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08724__A1 (.I(\u_cpu.rf_ram.memory[49][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06762__I1 (.I(\u_cpu.rf_ram.memory[49][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08726__A1 (.I(\u_cpu.rf_ram.memory[49][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06850__I1 (.I(\u_cpu.rf_ram.memory[49][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07654__A1 (.I(\u_cpu.rf_ram.memory[50][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06044__I2 (.I(\u_cpu.rf_ram.memory[50][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07656__A1 (.I(\u_cpu.rf_ram.memory[50][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06250__I2 (.I(\u_cpu.rf_ram.memory[50][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07659__A1 (.I(\u_cpu.rf_ram.memory[50][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06364__I2 (.I(\u_cpu.rf_ram.memory[50][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07661__A1 (.I(\u_cpu.rf_ram.memory[50][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06479__I2 (.I(\u_cpu.rf_ram.memory[50][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07663__A1 (.I(\u_cpu.rf_ram.memory[50][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06586__I2 (.I(\u_cpu.rf_ram.memory[50][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07665__A1 (.I(\u_cpu.rf_ram.memory[50][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06674__I2 (.I(\u_cpu.rf_ram.memory[50][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07667__A1 (.I(\u_cpu.rf_ram.memory[50][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06762__I2 (.I(\u_cpu.rf_ram.memory[50][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07669__A1 (.I(\u_cpu.rf_ram.memory[50][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06850__I2 (.I(\u_cpu.rf_ram.memory[50][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08272__A1 (.I(\u_cpu.rf_ram.memory[56][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06060__I0 (.I(\u_cpu.rf_ram.memory[56][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08276__A1 (.I(\u_cpu.rf_ram.memory[56][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06256__I0 (.I(\u_cpu.rf_ram.memory[56][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08281__A1 (.I(\u_cpu.rf_ram.memory[56][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06368__I0 (.I(\u_cpu.rf_ram.memory[56][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08285__A1 (.I(\u_cpu.rf_ram.memory[56][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06486__I0 (.I(\u_cpu.rf_ram.memory[56][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08289__A1 (.I(\u_cpu.rf_ram.memory[56][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06590__I0 (.I(\u_cpu.rf_ram.memory[56][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08293__A1 (.I(\u_cpu.rf_ram.memory[56][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06678__I0 (.I(\u_cpu.rf_ram.memory[56][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08297__A1 (.I(\u_cpu.rf_ram.memory[56][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06766__I0 (.I(\u_cpu.rf_ram.memory[56][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08301__A1 (.I(\u_cpu.rf_ram.memory[56][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06854__I0 (.I(\u_cpu.rf_ram.memory[56][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10922__A1 (.I(\u_cpu.rf_ram.memory[59][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06060__I3 (.I(\u_cpu.rf_ram.memory[59][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10924__A1 (.I(\u_cpu.rf_ram.memory[59][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06256__I3 (.I(\u_cpu.rf_ram.memory[59][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10927__A1 (.I(\u_cpu.rf_ram.memory[59][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06368__I3 (.I(\u_cpu.rf_ram.memory[59][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10929__A1 (.I(\u_cpu.rf_ram.memory[59][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06486__I3 (.I(\u_cpu.rf_ram.memory[59][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10931__A1 (.I(\u_cpu.rf_ram.memory[59][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06590__I3 (.I(\u_cpu.rf_ram.memory[59][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10933__A1 (.I(\u_cpu.rf_ram.memory[59][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06678__I3 (.I(\u_cpu.rf_ram.memory[59][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10935__A1 (.I(\u_cpu.rf_ram.memory[59][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06766__I3 (.I(\u_cpu.rf_ram.memory[59][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10937__A1 (.I(\u_cpu.rf_ram.memory[59][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06854__I3 (.I(\u_cpu.rf_ram.memory[59][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08172__A1 (.I(\u_cpu.rf_ram.memory[60][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06052__I0 (.I(\u_cpu.rf_ram.memory[60][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08174__A1 (.I(\u_cpu.rf_ram.memory[60][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06253__I0 (.I(\u_cpu.rf_ram.memory[60][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08123__A1 (.I(\u_cpu.rf_ram.memory[62][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06052__I2 (.I(\u_cpu.rf_ram.memory[62][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08125__A1 (.I(\u_cpu.rf_ram.memory[62][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06253__I2 (.I(\u_cpu.rf_ram.memory[62][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08128__A1 (.I(\u_cpu.rf_ram.memory[62][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06366__I2 (.I(\u_cpu.rf_ram.memory[62][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08130__A1 (.I(\u_cpu.rf_ram.memory[62][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06482__I2 (.I(\u_cpu.rf_ram.memory[62][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08132__A1 (.I(\u_cpu.rf_ram.memory[62][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06588__I2 (.I(\u_cpu.rf_ram.memory[62][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08134__A1 (.I(\u_cpu.rf_ram.memory[62][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06676__I2 (.I(\u_cpu.rf_ram.memory[62][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08136__A1 (.I(\u_cpu.rf_ram.memory[62][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06764__I2 (.I(\u_cpu.rf_ram.memory[62][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08138__A1 (.I(\u_cpu.rf_ram.memory[62][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06852__I2 (.I(\u_cpu.rf_ram.memory[62][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08108__A1 (.I(\u_cpu.rf_ram.memory[63][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06366__I3 (.I(\u_cpu.rf_ram.memory[63][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08110__A1 (.I(\u_cpu.rf_ram.memory[63][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06482__I3 (.I(\u_cpu.rf_ram.memory[63][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08112__A1 (.I(\u_cpu.rf_ram.memory[63][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06588__I3 (.I(\u_cpu.rf_ram.memory[63][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08118__A1 (.I(\u_cpu.rf_ram.memory[63][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06852__I3 (.I(\u_cpu.rf_ram.memory[63][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08061__A1 (.I(\u_cpu.rf_ram.memory[64][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06172__I0 (.I(\u_cpu.rf_ram.memory[64][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08063__A1 (.I(\u_cpu.rf_ram.memory[64][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06311__I0 (.I(\u_cpu.rf_ram.memory[64][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08066__A1 (.I(\u_cpu.rf_ram.memory[64][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06426__I0 (.I(\u_cpu.rf_ram.memory[64][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08068__A1 (.I(\u_cpu.rf_ram.memory[64][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06542__I0 (.I(\u_cpu.rf_ram.memory[64][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08070__A1 (.I(\u_cpu.rf_ram.memory[64][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06632__I0 (.I(\u_cpu.rf_ram.memory[64][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08072__A1 (.I(\u_cpu.rf_ram.memory[64][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06720__I0 (.I(\u_cpu.rf_ram.memory[64][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08074__A1 (.I(\u_cpu.rf_ram.memory[64][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06808__I0 (.I(\u_cpu.rf_ram.memory[64][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08076__A1 (.I(\u_cpu.rf_ram.memory[64][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06896__I0 (.I(\u_cpu.rf_ram.memory[64][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08047__A1 (.I(\u_cpu.rf_ram.memory[65][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06632__I1 (.I(\u_cpu.rf_ram.memory[65][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08050__A1 (.I(\u_cpu.rf_ram.memory[65][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06720__I1 (.I(\u_cpu.rf_ram.memory[65][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08053__A1 (.I(\u_cpu.rf_ram.memory[65][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06808__I1 (.I(\u_cpu.rf_ram.memory[65][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08056__A1 (.I(\u_cpu.rf_ram.memory[65][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06896__I1 (.I(\u_cpu.rf_ram.memory[65][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07972__A1 (.I(\u_cpu.rf_ram.memory[68][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06177__I0 (.I(\u_cpu.rf_ram.memory[68][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08584__A1 (.I(\u_cpu.rf_ram.memory[70][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06177__I2 (.I(\u_cpu.rf_ram.memory[70][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08586__A1 (.I(\u_cpu.rf_ram.memory[70][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06315__I2 (.I(\u_cpu.rf_ram.memory[70][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08589__A1 (.I(\u_cpu.rf_ram.memory[70][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06428__I2 (.I(\u_cpu.rf_ram.memory[70][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08591__A1 (.I(\u_cpu.rf_ram.memory[70][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06544__I2 (.I(\u_cpu.rf_ram.memory[70][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08593__A1 (.I(\u_cpu.rf_ram.memory[70][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06634__I2 (.I(\u_cpu.rf_ram.memory[70][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08595__A1 (.I(\u_cpu.rf_ram.memory[70][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06722__I2 (.I(\u_cpu.rf_ram.memory[70][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08597__A1 (.I(\u_cpu.rf_ram.memory[70][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06810__I2 (.I(\u_cpu.rf_ram.memory[70][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08599__A1 (.I(\u_cpu.rf_ram.memory[70][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06898__I2 (.I(\u_cpu.rf_ram.memory[70][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08557__A1 (.I(\u_cpu.rf_ram.memory[71][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06177__I3 (.I(\u_cpu.rf_ram.memory[71][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08560__A1 (.I(\u_cpu.rf_ram.memory[71][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06315__I3 (.I(\u_cpu.rf_ram.memory[71][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08564__A1 (.I(\u_cpu.rf_ram.memory[71][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06428__I3 (.I(\u_cpu.rf_ram.memory[71][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08567__A1 (.I(\u_cpu.rf_ram.memory[71][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06544__I3 (.I(\u_cpu.rf_ram.memory[71][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08570__A1 (.I(\u_cpu.rf_ram.memory[71][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06634__I3 (.I(\u_cpu.rf_ram.memory[71][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08573__A1 (.I(\u_cpu.rf_ram.memory[71][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06722__I3 (.I(\u_cpu.rf_ram.memory[71][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08576__A1 (.I(\u_cpu.rf_ram.memory[71][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06810__I3 (.I(\u_cpu.rf_ram.memory[71][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08579__A1 (.I(\u_cpu.rf_ram.memory[71][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06898__I3 (.I(\u_cpu.rf_ram.memory[71][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08516__A1 (.I(\u_cpu.rf_ram.memory[72][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06183__I0 (.I(\u_cpu.rf_ram.memory[72][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08518__A1 (.I(\u_cpu.rf_ram.memory[72][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06319__I0 (.I(\u_cpu.rf_ram.memory[72][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08521__A1 (.I(\u_cpu.rf_ram.memory[72][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06430__I0 (.I(\u_cpu.rf_ram.memory[72][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08523__A1 (.I(\u_cpu.rf_ram.memory[72][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06546__I0 (.I(\u_cpu.rf_ram.memory[72][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08525__A1 (.I(\u_cpu.rf_ram.memory[72][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06636__I0 (.I(\u_cpu.rf_ram.memory[72][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08527__A1 (.I(\u_cpu.rf_ram.memory[72][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06724__I0 (.I(\u_cpu.rf_ram.memory[72][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08529__A1 (.I(\u_cpu.rf_ram.memory[72][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06812__I0 (.I(\u_cpu.rf_ram.memory[72][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08531__A1 (.I(\u_cpu.rf_ram.memory[72][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06900__I0 (.I(\u_cpu.rf_ram.memory[72][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08536__A1 (.I(\u_cpu.rf_ram.memory[73][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06183__I1 (.I(\u_cpu.rf_ram.memory[73][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08538__A1 (.I(\u_cpu.rf_ram.memory[73][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06319__I1 (.I(\u_cpu.rf_ram.memory[73][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08541__A1 (.I(\u_cpu.rf_ram.memory[73][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06430__I1 (.I(\u_cpu.rf_ram.memory[73][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08543__A1 (.I(\u_cpu.rf_ram.memory[73][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06546__I1 (.I(\u_cpu.rf_ram.memory[73][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08545__A1 (.I(\u_cpu.rf_ram.memory[73][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06636__I1 (.I(\u_cpu.rf_ram.memory[73][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08547__A1 (.I(\u_cpu.rf_ram.memory[73][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06724__I1 (.I(\u_cpu.rf_ram.memory[73][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08549__A1 (.I(\u_cpu.rf_ram.memory[73][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06812__I1 (.I(\u_cpu.rf_ram.memory[73][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08551__A1 (.I(\u_cpu.rf_ram.memory[73][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06900__I1 (.I(\u_cpu.rf_ram.memory[73][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07884__A1 (.I(\u_cpu.rf_ram.memory[74][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06319__I2 (.I(\u_cpu.rf_ram.memory[74][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07891__A1 (.I(\u_cpu.rf_ram.memory[74][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06636__I2 (.I(\u_cpu.rf_ram.memory[74][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07906__A1 (.I(\u_cpu.rf_ram.memory[76][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06321__I0 (.I(\u_cpu.rf_ram.memory[76][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07919__A1 (.I(\u_cpu.rf_ram.memory[76][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06726__I0 (.I(\u_cpu.rf_ram.memory[76][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07409__A1 (.I(\u_cpu.rf_ram.memory[78][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06187__I2 (.I(\u_cpu.rf_ram.memory[78][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07411__A1 (.I(\u_cpu.rf_ram.memory[78][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06321__I2 (.I(\u_cpu.rf_ram.memory[78][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10745__A1 (.I(\u_cpu.rf_ram.memory[79][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06187__I3 (.I(\u_cpu.rf_ram.memory[79][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10748__A1 (.I(\u_cpu.rf_ram.memory[79][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06321__I3 (.I(\u_cpu.rf_ram.memory[79][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10752__A1 (.I(\u_cpu.rf_ram.memory[79][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06433__I3 (.I(\u_cpu.rf_ram.memory[79][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10758__A1 (.I(\u_cpu.rf_ram.memory[79][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06638__I3 (.I(\u_cpu.rf_ram.memory[79][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10764__A1 (.I(\u_cpu.rf_ram.memory[79][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06814__I3 (.I(\u_cpu.rf_ram.memory[79][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10767__A1 (.I(\u_cpu.rf_ram.memory[79][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06902__I3 (.I(\u_cpu.rf_ram.memory[79][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07386__A1 (.I(\u_cpu.rf_ram.memory[80][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06627__I0 (.I(\u_cpu.rf_ram.memory[80][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07186__A1 (.I(\u_cpu.rf_ram.memory[82][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06627__I2 (.I(\u_cpu.rf_ram.memory[82][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10835__A1 (.I(\u_cpu.rf_ram.memory[83][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06304__I3 (.I(\u_cpu.rf_ram.memory[83][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10846__A1 (.I(\u_cpu.rf_ram.memory[83][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06803__I3 (.I(\u_cpu.rf_ram.memory[83][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10848__A1 (.I(\u_cpu.rf_ram.memory[83][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06891__I3 (.I(\u_cpu.rf_ram.memory[83][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10902__A1 (.I(\u_cpu.rf_ram.memory[84][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06164__I0 (.I(\u_cpu.rf_ram.memory[84][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10904__A1 (.I(\u_cpu.rf_ram.memory[84][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06307__I0 (.I(\u_cpu.rf_ram.memory[84][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10907__A1 (.I(\u_cpu.rf_ram.memory[84][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06421__I0 (.I(\u_cpu.rf_ram.memory[84][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10909__A1 (.I(\u_cpu.rf_ram.memory[84][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06538__I0 (.I(\u_cpu.rf_ram.memory[84][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10913__A1 (.I(\u_cpu.rf_ram.memory[84][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06717__I0 (.I(\u_cpu.rf_ram.memory[84][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11008__A1 (.I(\u_cpu.rf_ram.memory[86][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06164__I2 (.I(\u_cpu.rf_ram.memory[86][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11010__A1 (.I(\u_cpu.rf_ram.memory[86][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06307__I2 (.I(\u_cpu.rf_ram.memory[86][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11015__A1 (.I(\u_cpu.rf_ram.memory[86][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06538__I2 (.I(\u_cpu.rf_ram.memory[86][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11017__A1 (.I(\u_cpu.rf_ram.memory[86][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06629__I2 (.I(\u_cpu.rf_ram.memory[86][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11021__A1 (.I(\u_cpu.rf_ram.memory[86][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06805__I2 (.I(\u_cpu.rf_ram.memory[86][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11023__A1 (.I(\u_cpu.rf_ram.memory[86][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06893__I2 (.I(\u_cpu.rf_ram.memory[86][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11061__A1 (.I(\u_cpu.rf_ram.memory[87][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06805__I3 (.I(\u_cpu.rf_ram.memory[87][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11063__A1 (.I(\u_cpu.rf_ram.memory[87][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06893__I3 (.I(\u_cpu.rf_ram.memory[87][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11073__A1 (.I(\u_cpu.rf_ram.memory[88][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06415__I0 (.I(\u_cpu.rf_ram.memory[88][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11075__A1 (.I(\u_cpu.rf_ram.memory[88][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06531__I0 (.I(\u_cpu.rf_ram.memory[88][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11077__A1 (.I(\u_cpu.rf_ram.memory[88][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06625__I0 (.I(\u_cpu.rf_ram.memory[88][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11079__A1 (.I(\u_cpu.rf_ram.memory[88][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06713__I0 (.I(\u_cpu.rf_ram.memory[88][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11081__A1 (.I(\u_cpu.rf_ram.memory[88][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06801__I0 (.I(\u_cpu.rf_ram.memory[88][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11083__A1 (.I(\u_cpu.rf_ram.memory[88][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06889__I0 (.I(\u_cpu.rf_ram.memory[88][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11282__A1 (.I(\u_cpu.rf_ram.memory[89][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06625__I1 (.I(\u_cpu.rf_ram.memory[89][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11284__A1 (.I(\u_cpu.rf_ram.memory[89][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06713__I1 (.I(\u_cpu.rf_ram.memory[89][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11288__A1 (.I(\u_cpu.rf_ram.memory[89][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06889__I1 (.I(\u_cpu.rf_ram.memory[89][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09366__I1 (.I(\u_cpu.rf_ram.memory[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05961__I0 (.I(\u_cpu.rf_ram.memory[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09171__A1 (.I(\u_cpu.rf_ram.memory[90][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06152__I2 (.I(\u_cpu.rf_ram.memory[90][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09174__A1 (.I(\u_cpu.rf_ram.memory[90][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06302__I2 (.I(\u_cpu.rf_ram.memory[90][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09184__A1 (.I(\u_cpu.rf_ram.memory[90][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06625__I2 (.I(\u_cpu.rf_ram.memory[90][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09150__A1 (.I(\u_cpu.rf_ram.memory[91][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06152__I3 (.I(\u_cpu.rf_ram.memory[91][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09152__A1 (.I(\u_cpu.rf_ram.memory[91][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06302__I3 (.I(\u_cpu.rf_ram.memory[91][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09155__A1 (.I(\u_cpu.rf_ram.memory[91][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06415__I3 (.I(\u_cpu.rf_ram.memory[91][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09157__A1 (.I(\u_cpu.rf_ram.memory[91][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06531__I3 (.I(\u_cpu.rf_ram.memory[91][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09159__A1 (.I(\u_cpu.rf_ram.memory[91][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06625__I3 (.I(\u_cpu.rf_ram.memory[91][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09161__A1 (.I(\u_cpu.rf_ram.memory[91][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06713__I3 (.I(\u_cpu.rf_ram.memory[91][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09163__A1 (.I(\u_cpu.rf_ram.memory[91][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06801__I3 (.I(\u_cpu.rf_ram.memory[91][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09218__A1 (.I(\u_cpu.rf_ram.memory[92][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06147__I0 (.I(\u_cpu.rf_ram.memory[92][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09220__A1 (.I(\u_cpu.rf_ram.memory[92][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06300__I0 (.I(\u_cpu.rf_ram.memory[92][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09223__A1 (.I(\u_cpu.rf_ram.memory[92][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06412__I0 (.I(\u_cpu.rf_ram.memory[92][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09225__A1 (.I(\u_cpu.rf_ram.memory[92][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06529__I0 (.I(\u_cpu.rf_ram.memory[92][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09229__A1 (.I(\u_cpu.rf_ram.memory[92][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06711__I0 (.I(\u_cpu.rf_ram.memory[92][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10514__A1 (.I(\u_cpu.rf_ram.memory[94][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06147__I2 (.I(\u_cpu.rf_ram.memory[94][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10516__A1 (.I(\u_cpu.rf_ram.memory[94][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06300__I2 (.I(\u_cpu.rf_ram.memory[94][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10519__A1 (.I(\u_cpu.rf_ram.memory[94][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06412__I2 (.I(\u_cpu.rf_ram.memory[94][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10521__A1 (.I(\u_cpu.rf_ram.memory[94][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06529__I2 (.I(\u_cpu.rf_ram.memory[94][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10523__A1 (.I(\u_cpu.rf_ram.memory[94][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06623__I2 (.I(\u_cpu.rf_ram.memory[94][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10525__A1 (.I(\u_cpu.rf_ram.memory[94][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06711__I2 (.I(\u_cpu.rf_ram.memory[94][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10527__A1 (.I(\u_cpu.rf_ram.memory[94][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06799__I2 (.I(\u_cpu.rf_ram.memory[94][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10529__A1 (.I(\u_cpu.rf_ram.memory[94][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06887__I2 (.I(\u_cpu.rf_ram.memory[94][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10543__A1 (.I(\u_cpu.rf_ram.memory[95][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06623__I3 (.I(\u_cpu.rf_ram.memory[95][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10545__A1 (.I(\u_cpu.rf_ram.memory[95][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06711__I3 (.I(\u_cpu.rf_ram.memory[95][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10547__A1 (.I(\u_cpu.rf_ram.memory[95][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06799__I3 (.I(\u_cpu.rf_ram.memory[95][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10549__A1 (.I(\u_cpu.rf_ram.memory[95][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06887__I3 (.I(\u_cpu.rf_ram.memory[95][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10559__A1 (.I(\u_cpu.rf_ram.memory[96][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06396__I0 (.I(\u_cpu.rf_ram.memory[96][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10561__A1 (.I(\u_cpu.rf_ram.memory[96][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06512__I0 (.I(\u_cpu.rf_ram.memory[96][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10563__A1 (.I(\u_cpu.rf_ram.memory[96][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06610__I0 (.I(\u_cpu.rf_ram.memory[96][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10565__A1 (.I(\u_cpu.rf_ram.memory[96][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06698__I0 (.I(\u_cpu.rf_ram.memory[96][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10567__A1 (.I(\u_cpu.rf_ram.memory[96][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06786__I0 (.I(\u_cpu.rf_ram.memory[96][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11233__A1 (.I(\u_cpu.rf_ram.memory[98][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06113__I2 (.I(\u_cpu.rf_ram.memory[98][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11235__A1 (.I(\u_cpu.rf_ram.memory[98][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06282__I2 (.I(\u_cpu.rf_ram.memory[98][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11238__A1 (.I(\u_cpu.rf_ram.memory[98][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06396__I2 (.I(\u_cpu.rf_ram.memory[98][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11240__A1 (.I(\u_cpu.rf_ram.memory[98][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06512__I2 (.I(\u_cpu.rf_ram.memory[98][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11242__A1 (.I(\u_cpu.rf_ram.memory[98][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06610__I2 (.I(\u_cpu.rf_ram.memory[98][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10731__A1 (.I(\u_cpu.rf_ram.memory[99][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06512__I3 (.I(\u_cpu.rf_ram.memory[99][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08389__I1 (.I(\u_cpu.rf_ram.memory[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06223__I1 (.I(\u_cpu.rf_ram.memory[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08392__I1 (.I(\u_cpu.rf_ram.memory[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06339__I1 (.I(\u_cpu.rf_ram.memory[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08395__I1 (.I(\u_cpu.rf_ram.memory[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06452__I1 (.I(\u_cpu.rf_ram.memory[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08407__I1 (.I(\u_cpu.rf_ram.memory[9][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06830__I1 (.I(\u_cpu.rf_ram.memory[9][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07144__I (.I(\u_cpu.rf_ram_if.genblk1.wtrig0_r ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07130__I (.I(\u_cpu.rf_ram_if.genblk1.wtrig0_r ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07127__A1 (.I(\u_cpu.rf_ram_if.genblk1.wtrig0_r ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07126__B (.I(\u_cpu.rf_ram_if.genblk1.wtrig0_r ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12695__D (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11315__A3 (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07145__B1 (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05764__B (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05756__A2 (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12685__D (.I(\u_cpu.rf_ram_if.wdata0_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07317__I0 (.I(\u_cpu.rf_ram_if.wdata0_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07170__A2 (.I(\u_cpu.rf_ram_if.wdata0_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12687__D (.I(\u_cpu.rf_ram_if.wdata0_r[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07325__I0 (.I(\u_cpu.rf_ram_if.wdata0_r[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07183__A2 (.I(\u_cpu.rf_ram_if.wdata0_r[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12698__D (.I(\u_cpu.rf_ram_if.wdata1_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07317__I1 (.I(\u_cpu.rf_ram_if.wdata1_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07169__A2 (.I(\u_cpu.rf_ram_if.wdata1_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12700__D (.I(\u_cpu.rf_ram_if.wdata1_r[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07325__I1 (.I(\u_cpu.rf_ram_if.wdata1_r[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07182__A2 (.I(\u_cpu.rf_ram_if.wdata1_r[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12703__D (.I(\u_cpu.rf_ram_if.wdata1_r[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07337__I0 (.I(\u_cpu.rf_ram_if.wdata1_r[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07200__A2 (.I(\u_cpu.rf_ram_if.wdata1_r[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout35_I (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[38]_D  (.I(\u_scanchain_local.module_data_in[37] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.out_flop_D  (.I(\u_scanchain_local.module_data_in[69] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10283__A1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10280__B (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09136__A1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07689__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05783__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[0]_D  (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout565_I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output7_I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07711__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[2]_D  (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09527__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09740__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07694__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[19]_CLK  (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[18]_CLK  (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[24]_CLK  (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[20]_CLK  (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[21]_CLK  (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout10_I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[17]_CLK  (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[15]_CLK  (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[16]_CLK  (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[14]_CLK  (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[22]_CLK  (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[29]_CLK  (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[26]_CLK  (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[27]_CLK  (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout12_I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout13_I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout9_I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout11_I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[7]_CLK  (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[6]_CLK  (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[2]_CLK  (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[5]_CLK  (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[4]_CLK  (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[34]_CLK  (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[35]_CLK  (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[32]_CLK  (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[8]_CLK  (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout15_I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[28]_CLK  (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[33]_CLK  (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[3]_CLK  (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[31]_CLK  (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[30]_CLK  (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout16_I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout17_I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout18_I (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout14_I (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[40]_CLK  (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[38]_CLK  (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[0]_CLK  (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[1]_CLK  (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[39]_CLK  (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[62]_CLK  (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[60]_CLK  (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[66]_CLK  (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[65]_CLK  (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[67]_CLK  (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[64]_CLK  (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[61]_CLK  (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout22_I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout23_I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[36]_CLK  (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[63]_CLK  (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[37]_CLK  (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout24_I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout20_I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout21_I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[47]_CLK  (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[48]_CLK  (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[50]_CLK  (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.out_flop_CLKN  (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[46]_CLK  (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[45]_CLK  (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[44]_CLK  (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[43]_CLK  (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[69]_CLK  (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[68]_CLK  (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[49]_CLK  (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout26_I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout29_I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout30_I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[59]_CLK  (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[57]_CLK  (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout31_I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout27_I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout28_I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout32_I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout25_I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout33_I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.output_buffers[3]_I  (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout34_I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout19_I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12461__CLK (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12459__CLK (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12458__CLK (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12500__CLK (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12499__CLK (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12502__CLK (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12501__CLK (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12494__CLK (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12486__CLK (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12497__CLK (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12489__CLK (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12484__CLK (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12483__CLK (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12482__CLK (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout40_I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout41_I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout38_I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout39_I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout42_I (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12462__CLK (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout37_I (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12467__CLK (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout44_I (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12460__CLK (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12457__CLK (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12456__CLK (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout47_I (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12487__CLK (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12481__CLK (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12480__CLK (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12463__CLK (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout46_I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout48_I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout45_I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout49_I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout43_I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12621__CLK (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12620__CLK (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12614__CLK (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12613__CLK (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12612__CLK (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12626__CLK (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12630__CLK (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12629__CLK (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12628__CLK (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12622__CLK (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout53_I (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout54_I (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout51_I (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout52_I (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11357__CLK (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11356__CLK (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12617__CLK (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12616__CLK (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12615__CLK (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11665__CLK (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout56_I (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout57_I (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout59_I (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout60_I (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout58_I (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout61_I (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout55_I (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12651__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12650__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11361__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout63_I (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout64_I (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11477__CLK (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11350__CLK (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11348__CLK (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12640__CLK (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11354__CLK (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11360__CLK (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11359__CLK (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11355__CLK (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11331__CLK (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11330__CLK (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11352__CLK (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11351__CLK (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11349__CLK (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11347__CLK (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout68_I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout69_I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11666__CLK (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout67_I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout70_I (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout65_I (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout66_I (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout71_I (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout62_I (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12404__CLK (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12403__CLK (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12377__CLK (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12375__CLK (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12374__CLK (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12405__CLK (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout74_I (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12402__CLK (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12401__CLK (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12381__CLK (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12445__CLK (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12444__CLK (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12443__CLK (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12442__CLK (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12379__CLK (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12300__CLK (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12258__CLK (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12378__CLK (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12376__CLK (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12299__CLK (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12257__CLK (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12412__CLK (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12409__CLK (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12408__CLK (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout81_I (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout82_I (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout79_I (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout80_I (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout83_I (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout78_I (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12454__CLK (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12439__CLK (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12438__CLK (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12453__CLK (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12437__CLK (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout87_I (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout88_I (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout85_I (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout86_I (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12413__CLK (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12411__CLK (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12410__CLK (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12301__CLK (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12259__CLK (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11326__CLK (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout90_I (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout89_I (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout91_I (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout84_I (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12256__CLK (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12253__CLK (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12654__CLK (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12295__CLK (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12252__CLK (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12678__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12677__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11337__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout93_I (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout94_I (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12681__CLK (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12296__CLK (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12254__CLK (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout95_I (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout96_I (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11494__CLK (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11353__CLK (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11346__CLK (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11336__CLK (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11335__CLK (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11502__CLK (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11495__CLK (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11487__CLK (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11670__CLK (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout98_I (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout99_I (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12682__CLK (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout97_I (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11616__CLK (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11615__CLK (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11621__CLK (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11620__CLK (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11325__CLK (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout101_I (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout102_I (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11493__CLK (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11492__CLK (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11488__CLK (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout103_I (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout104_I (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout105_I (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout106_I (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout100_I (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout108_I (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout73_I (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11474__CLK (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11569__CLK (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11567__CLK (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11372__CLK (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11370__CLK (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12642__CLK (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12353__CLK (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12345__CLK (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11364__CLK (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11362__CLK (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12644__CLK (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout112_I (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout110_I (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout111_I (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11568__CLK (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11371__CLK (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11363__CLK (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11667__CLK (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11571__CLK (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12643__CLK (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout114_I (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout113_I (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12546__CLK (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12115__CLK (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12355__CLK (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12347__CLK (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12116__CLK (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout117_I (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout118_I (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12547__CLK (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout116_I (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout119_I (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout115_I (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11475__CLK (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11365__CLK (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11664__CLK (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11478__CLK (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11374__CLK (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11366__CLK (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11668__CLK (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11572__CLK (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11479__CLK (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11375__CLK (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout122_I (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout123_I (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12645__CLK (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout121_I (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12113__CLK (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12106__CLK (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12105__CLK (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12357__CLK (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12349__CLK (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11727__CLK (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12549__CLK (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12358__CLK (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12118__CLK (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12110__CLK (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout127_I (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout128_I (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout125_I (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout126_I (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout129_I (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout124_I (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout130_I (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout120_I (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11731__CLK (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout131_I (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12647__CLK (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11574__CLK (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11481__CLK (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11377__CLK (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11369__CLK (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12649__CLK (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11573__CLK (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11376__CLK (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11368__CLK (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12120__CLK (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12112__CLK (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11775__CLK (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout135_I (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout136_I (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout137_I (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout138_I (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout133_I (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout134_I (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11741__CLK (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12698__CLK (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12697__CLK (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12685__CLK (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11496__CLK (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout140_I (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout141_I (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12648__CLK (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11669__CLK (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11480__CLK (.I(net142));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11780__CLK (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11742__CLK (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11733__CLK (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout143_I (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout144_I (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout145_I (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout146_I (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout142_I (.I(net147));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout147_I (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout139_I (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11776__CLK (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11825__CLK (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11824__CLK (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11737__CLK (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11736__CLK (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11778__CLK (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11827__CLK (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11826__CLK (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11739__CLK (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11738__CLK (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout152_I (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout153_I (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout154_I (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout151_I (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout155_I (.I(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout148_I (.I(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout156_I (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout132_I (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout157_I (.I(net158));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout109_I (.I(net158));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12563__CLK (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12562__CLK (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12662__CLK (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12661__CLK (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12660__CLK (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12659__CLK (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12658__CLK (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12436__CLK (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12435__CLK (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12433__CLK (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12508__CLK (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12566__CLK (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12565__CLK (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12561__CLK (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12560__CLK (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12567__CLK (.I(net163));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout162_I (.I(net163));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12507__CLK (.I(net163));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12506__CLK (.I(net163));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout163_I (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout160_I (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout161_I (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12338__CLK (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12337__CLK (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12336__CLK (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout165_I (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout166_I (.I(net167));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12510__CLK (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12505__CLK (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12581__CLK (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12577__CLK (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12576__CLK (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12509__CLK (.I(net170));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11343__CLK (.I(net170));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11327__CLK (.I(net170));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout168_I (.I(net170));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout169_I (.I(net170));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout170_I (.I(net172));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout171_I (.I(net172));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12578__CLK (.I(net172));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout167_I (.I(net172));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout172_I (.I(net173));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout164_I (.I(net173));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11625__CLK (.I(net176));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11381__CLK (.I(net176));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11380__CLK (.I(net176));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout174_I (.I(net176));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout175_I (.I(net176));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12474__CLK (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11662__CLK (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11659__CLK (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11389__CLK (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout181_I (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout182_I (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout179_I (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout180_I (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout183_I (.I(net184));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout176_I (.I(net184));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout177_I (.I(net184));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11623__CLK (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12504__CLK (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11382__CLK (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11323__CLK (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11322__CLK (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11378__CLK (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11339__CLK (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11338__CLK (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout185_I (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout186_I (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11660__CLK (.I(net188));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11388__CLK (.I(net188));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11644__CLK (.I(net188));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11641__CLK (.I(net188));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11640__CLK (.I(net188));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11390__CLK (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11646__CLK (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11645__CLK (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11643__CLK (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11642__CLK (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout189_I (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout190_I (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11661__CLK (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout188_I (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout191_I (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout187_I (.I(net192));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout192_I (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout184_I (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12514__CLK (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12389__CLK (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12382__CLK (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12388__CLK (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout195_I (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12587__CLK (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12397__CLK (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12390__CLK (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12572__CLK (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12571__CLK (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout201_I (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout196_I (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout197_I (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12575__CLK (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12518__CLK (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12517__CLK (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12513__CLK (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12512__CLK (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12585__CLK (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12584__CLK (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11344__CLK (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout205_I (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout206_I (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout207_I (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout203_I (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout204_I (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout208_I (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout202_I (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12368__CLK (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12367__CLK (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12366__CLK (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12365__CLK (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12364__CLK (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout210_I (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12555__CLK (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12363__CLK (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12362__CLK (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12361__CLK (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12558__CLK (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12557__CLK (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12554__CLK (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12553__CLK (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12552__CLK (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12559__CLK (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout212_I (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12556__CLK (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout211_I (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11402__CLK (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11385__CLK (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11384__CLK (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11345__CLK (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11329__CLK (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout217_I (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout218_I (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout215_I (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout216_I (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11387__CLK (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11386__CLK (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11654__CLK (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11653__CLK (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11652__CLK (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11406__CLK (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11405__CLK (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11404__CLK (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11392__CLK (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout220_I (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout221_I (.I(net223));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout222_I (.I(net223));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout219_I (.I(net223));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11415__CLK (.I(net224));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11411__CLK (.I(net224));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11410__CLK (.I(net224));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11409__CLK (.I(net224));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11408__CLK (.I(net224));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11412__CLK (.I(net226));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11465__CLK (.I(net226));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11464__CLK (.I(net226));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11463__CLK (.I(net226));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11414__CLK (.I(net226));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout226_I (.I(net228));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout227_I (.I(net228));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout224_I (.I(net228));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout225_I (.I(net228));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout228_I (.I(net229));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout223_I (.I(net229));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout230_I (.I(net231));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout194_I (.I(net231));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12699__CLK (.I(net232));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12687__CLK (.I(net232));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12686__CLK (.I(net232));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12684__CLK (.I(net232));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12475__CLK (.I(net232));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12690__CLK (.I(net234));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12689__CLK (.I(net234));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12688__CLK (.I(net234));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11538__CLK (.I(net234));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12476__CLK (.I(net234));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12703__CLK (.I(net235));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout234_I (.I(net235));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout232_I (.I(net235));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout233_I (.I(net235));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11609__CLK (.I(net236));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11925__CLK (.I(net236));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11781__CLK (.I(net236));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11608__CLK (.I(net236));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11607__CLK (.I(net236));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11613__CLK (.I(net238));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11612__CLK (.I(net238));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11611__CLK (.I(net238));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout236_I (.I(net238));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout237_I (.I(net238));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12704__CLK (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11614__CLK (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout238_I (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout239_I (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout235_I (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12473__CLK (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12472__CLK (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11554__CLK (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11553__CLK (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11537__CLK (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12479__CLK (.I(net242));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11555__CLK (.I(net242));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11539__CLK (.I(net242));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11605__CLK (.I(net243));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11604__CLK (.I(net243));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11603__CLK (.I(net243));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11602__CLK (.I(net243));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11601__CLK (.I(net243));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11593__CLK (.I(net244));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout243_I (.I(net244));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11606__CLK (.I(net244));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11600__CLK (.I(net244));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11599__CLK (.I(net244));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11594__CLK (.I(net246));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout245_I (.I(net246));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout241_I (.I(net246));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout242_I (.I(net246));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout246_I (.I(net247));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout240_I (.I(net247));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11586__CLK (.I(net248));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11585__CLK (.I(net248));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout247_I (.I(net248));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11557__CLK (.I(net249));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11556__CLK (.I(net249));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11541__CLK (.I(net249));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11540__CLK (.I(net249));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11393__CLK (.I(net249));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11558__CLK (.I(net250));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11551__CLK (.I(net250));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11542__CLK (.I(net250));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11536__CLK (.I(net250));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11535__CLK (.I(net250));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11596__CLK (.I(net251));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11595__CLK (.I(net251));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11587__CLK (.I(net251));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11598__CLK (.I(net251));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11597__CLK (.I(net251));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout252_I (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11747__CLK (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11590__CLK (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11589__CLK (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11552__CLK (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11750__CLK (.I(net254));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout253_I (.I(net254));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11980__CLK (.I(net254));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout251_I (.I(net254));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout254_I (.I(net255));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout249_I (.I(net255));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout250_I (.I(net255));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12674__CLK (.I(net256));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11749__CLK (.I(net256));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11748__CLK (.I(net256));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11743__CLK (.I(net256));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11543__CLK (.I(net256));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12693__CLK (.I(net257));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11995__CLK (.I(net257));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11991__CLK (.I(net257));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11559__CLK (.I(net257));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout256_I (.I(net257));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11561__CLK (.I(net258));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11560__CLK (.I(net258));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11547__CLK (.I(net258));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11546__CLK (.I(net258));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11545__CLK (.I(net258));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11994__CLK (.I(net259));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11993__CLK (.I(net259));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11992__CLK (.I(net259));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11562__CLK (.I(net259));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout258_I (.I(net259));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12241__CLK (.I(net260));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout259_I (.I(net260));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12695__CLK (.I(net260));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout257_I (.I(net260));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout260_I (.I(net261));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11550__CLK (.I(net261));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11544__CLK (.I(net261));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout261_I (.I(net262));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout255_I (.I(net262));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12235__CLK (.I(net263));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12234__CLK (.I(net263));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11990__CLK (.I(net263));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11989__CLK (.I(net263));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11975__CLK (.I(net263));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12420__CLK (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12418__CLK (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12236__CLK (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout263_I (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout264_I (.I(net265));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11979__CLK (.I(net265));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11978__CLK (.I(net265));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11977__CLK (.I(net265));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11976__CLK (.I(net265));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout265_I (.I(net266));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout262_I (.I(net266));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout266_I (.I(net267));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout248_I (.I(net267));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout267_I (.I(net268));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout231_I (.I(net268));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout268_I (.I(net269));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout158_I (.I(net269));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12531__CLK (.I(net271));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12056__CLK (.I(net271));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12049__CLK (.I(net271));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12055__CLK (.I(net271));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout270_I (.I(net271));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12596__CLK (.I(net274));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12595__CLK (.I(net274));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12251__CLK (.I(net274));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12244__CLK (.I(net274));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout273_I (.I(net274));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout274_I (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12532__CLK (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout271_I (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12529__CLK (.I(net276));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12528__CLK (.I(net276));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12534__CLK (.I(net276));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12533__CLK (.I(net276));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12530__CLK (.I(net276));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12538__CLK (.I(net279));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout278_I (.I(net279));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12598__CLK (.I(net279));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12597__CLK (.I(net279));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12594__CLK (.I(net279));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout279_I (.I(net280));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout276_I (.I(net280));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout277_I (.I(net280));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout280_I (.I(net281));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout275_I (.I(net281));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12070__CLK (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12066__CLK (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12069__CLK (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12068__CLK (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12067__CLK (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12072__CLK (.I(net284));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12065__CLK (.I(net284));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12037__CLK (.I(net284));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12036__CLK (.I(net284));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout283_I (.I(net284));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12062__CLK (.I(net285));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12040__CLK (.I(net285));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12039__CLK (.I(net285));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12038__CLK (.I(net285));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout284_I (.I(net285));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11677__CLK (.I(net286));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12670__CLK (.I(net286));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12669__CLK (.I(net286));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12668__CLK (.I(net286));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12666__CLK (.I(net286));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12672__CLK (.I(net288));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12671__CLK (.I(net288));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11676__CLK (.I(net288));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout286_I (.I(net288));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout287_I (.I(net288));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12673__CLK (.I(net289));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout288_I (.I(net289));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12064__CLK (.I(net289));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout285_I (.I(net289));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout289_I (.I(net290));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout281_I (.I(net290));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11422__CLK (.I(net291));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11419__CLK (.I(net291));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12543__CLK (.I(net291));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11425__CLK (.I(net291));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11418__CLK (.I(net291));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11400__CLK (.I(net293));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11399__CLK (.I(net293));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12541__CLK (.I(net293));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12540__CLK (.I(net293));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12539__CLK (.I(net293));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11401__CLK (.I(net294));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout293_I (.I(net294));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout291_I (.I(net294));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout292_I (.I(net294));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11504__CLK (.I(net295));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11503__CLK (.I(net295));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11443__CLK (.I(net295));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11442__CLK (.I(net295));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11395__CLK (.I(net295));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout296_I (.I(net297));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11462__CLK (.I(net297));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11421__CLK (.I(net297));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11420__CLK (.I(net297));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11394__CLK (.I(net297));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout295_I (.I(net298));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout297_I (.I(net298));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout294_I (.I(net298));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11397__CLK (.I(net299));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11686__CLK (.I(net299));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11678__CLK (.I(net299));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11449__CLK (.I(net299));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11448__CLK (.I(net299));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11684__CLK (.I(net300));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11447__CLK (.I(net300));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11467__CLK (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11466__CLK (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11510__CLK (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11509__CLK (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11398__CLK (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11469__CLK (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11468__CLK (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11507__CLK (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11505__CLK (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11396__CLK (.I(net302));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11508__CLK (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout302_I (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11473__CLK (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout301_I (.I(net303));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout303_I (.I(net304));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout299_I (.I(net304));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout300_I (.I(net304));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout304_I (.I(net305));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout298_I (.I(net305));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12153__CLK (.I(net310));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12077__CLK (.I(net310));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12073__CLK (.I(net310));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12159__CLK (.I(net310));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout309_I (.I(net310));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12160__CLK (.I(net311));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout310_I (.I(net311));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout307_I (.I(net311));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout308_I (.I(net311));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout313_I (.I(net314));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11679__CLK (.I(net314));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11673__CLK (.I(net314));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11672__CLK (.I(net314));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11671__CLK (.I(net314));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout312_I (.I(net315));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout314_I (.I(net315));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout311_I (.I(net315));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12219__CLK (.I(net318));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12213__CLK (.I(net318));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12212__CLK (.I(net318));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12076__CLK (.I(net318));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12075__CLK (.I(net318));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11512__CLK (.I(net319));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12079__CLK (.I(net319));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12078__CLK (.I(net319));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12034__CLK (.I(net319));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12033__CLK (.I(net319));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11514__CLK (.I(net320));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11513__CLK (.I(net320));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11511__CLK (.I(net320));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12028__CLK (.I(net320));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout319_I (.I(net320));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11518__CLK (.I(net321));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11515__CLK (.I(net321));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout320_I (.I(net322));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout321_I (.I(net322));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout317_I (.I(net322));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout318_I (.I(net322));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout322_I (.I(net323));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout315_I (.I(net323));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11440__CLK (.I(net324));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11437__CLK (.I(net324));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11683__CLK (.I(net324));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11682__CLK (.I(net324));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11681__CLK (.I(net324));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11441__CLK (.I(net325));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout324_I (.I(net325));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11675__CLK (.I(net325));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11674__CLK (.I(net325));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11445__CLK (.I(net325));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11426__CLK (.I(net326));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11506__CLK (.I(net326));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11446__CLK (.I(net326));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11444__CLK (.I(net326));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11433__CLK (.I(net326));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11457__CLK (.I(net327));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11436__CLK (.I(net327));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11434__CLK (.I(net327));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11429__CLK (.I(net327));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout326_I (.I(net328));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout327_I (.I(net328));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout325_I (.I(net328));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11719__CLK (.I(net332));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout331_I (.I(net332));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout329_I (.I(net332));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout330_I (.I(net332));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11428__CLK (.I(net333));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11934__CLK (.I(net333));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11932__CLK (.I(net333));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11928__CLK (.I(net333));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11451__CLK (.I(net333));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout333_I (.I(net334));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11454__CLK (.I(net334));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11453__CLK (.I(net334));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11450__CLK (.I(net334));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11435__CLK (.I(net334));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11452__CLK (.I(net335));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout334_I (.I(net335));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout332_I (.I(net335));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout335_I (.I(net336));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout328_I (.I(net336));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout337_I (.I(net338));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout306_I (.I(net338));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11581__CLK (.I(net339));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11549__CLK (.I(net339));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11548__CLK (.I(net339));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12527__CLK (.I(net339));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12526__CLK (.I(net339));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11580__CLK (.I(net340));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11576__CLK (.I(net340));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11575__CLK (.I(net340));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11582__CLK (.I(net340));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout339_I (.I(net340));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12239__CLK (.I(net341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12238__CLK (.I(net341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11563__CLK (.I(net341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11566__CLK (.I(net341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11565__CLK (.I(net341));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12372__CLK (.I(net343));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12371__CLK (.I(net343));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12224__CLK (.I(net343));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12223__CLK (.I(net343));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11564__CLK (.I(net343));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12373__CLK (.I(net344));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout343_I (.I(net344));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout341_I (.I(net344));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout342_I (.I(net344));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout344_I (.I(net345));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12525__CLK (.I(net345));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout340_I (.I(net345));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11790__CLK (.I(net347));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11577__CLK (.I(net347));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11806__CLK (.I(net347));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11805__CLK (.I(net347));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11470__CLK (.I(net347));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout347_I (.I(net349));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout348_I (.I(net349));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11578__CLK (.I(net349));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout346_I (.I(net349));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12221__CLK (.I(net350));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11787__CLK (.I(net350));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11786__CLK (.I(net350));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11785__CLK (.I(net350));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11579__CLK (.I(net350));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12210__CLK (.I(net352));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11794__CLK (.I(net352));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11793__CLK (.I(net352));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11784__CLK (.I(net352));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11783__CLK (.I(net352));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12706__CLK (.I(net353));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12705__CLK (.I(net353));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12220__CLK (.I(net353));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12211__CLK (.I(net353));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout352_I (.I(net354));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout353_I (.I(net354));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout350_I (.I(net354));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout351_I (.I(net354));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout354_I (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout349_I (.I(net355));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout355_I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout345_I (.I(net356));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12416__CLK (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12424__CLK (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12423__CLK (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12419__CLK (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12417__CLK (.I(net357));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout358_I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12370__CLK (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12237__CLK (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12233__CLK (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12225__CLK (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12228__CLK (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12227__CLK (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12608__CLK (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12232__CLK (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12202__CLK (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout360_I (.I(net362));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout361_I (.I(net362));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12226__CLK (.I(net362));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12204__CLK (.I(net362));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12174__CLK (.I(net363));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12430__CLK (.I(net363));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12429__CLK (.I(net363));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12425__CLK (.I(net363));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12422__CLK (.I(net363));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout363_I (.I(net365));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout364_I (.I(net365));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout362_I (.I(net365));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout365_I (.I(net366));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout357_I (.I(net366));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout359_I (.I(net366));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout366_I (.I(net367));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout356_I (.I(net367));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11801__CLK (.I(net368));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11798__CLK (.I(net368));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11799__CLK (.I(net368));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11432__CLK (.I(net368));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11431__CLK (.I(net368));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11814__CLK (.I(net370));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11807__CLK (.I(net370));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11456__CLK (.I(net370));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11455__CLK (.I(net370));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11430__CLK (.I(net370));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout370_I (.I(net372));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout371_I (.I(net372));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout368_I (.I(net372));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout369_I (.I(net372));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12602__CLK (.I(net373));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12209__CLK (.I(net373));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11795__CLK (.I(net373));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11792__CLK (.I(net373));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11791__CLK (.I(net373));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12601__CLK (.I(net374));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11796__CLK (.I(net374));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11788__CLK (.I(net374));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12603__CLK (.I(net374));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout373_I (.I(net374));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout374_I (.I(net375));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout372_I (.I(net375));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11486__CLK (.I(net376));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11812__CLK (.I(net376));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11811__CLK (.I(net376));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11808__CLK (.I(net376));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11485__CLK (.I(net376));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12605__CLK (.I(net378));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12604__CLK (.I(net378));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12600__CLK (.I(net378));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11484__CLK (.I(net378));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11483__CLK (.I(net378));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12048__CLK (.I(net379));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12020__CLK (.I(net379));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11482__CLK (.I(net379));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12696__CLK (.I(net379));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12694__CLK (.I(net379));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12609__CLK (.I(net380));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout379_I (.I(net380));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12607__CLK (.I(net380));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout378_I (.I(net380));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout380_I (.I(net381));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout376_I (.I(net381));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout377_I (.I(net381));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout381_I (.I(net382));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout375_I (.I(net382));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12206__CLK (.I(net383));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12170__CLK (.I(net383));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12406__CLK (.I(net383));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12242__CLK (.I(net383));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12231__CLK (.I(net383));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout383_I (.I(net384));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12208__CLK (.I(net384));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12205__CLK (.I(net384));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12203__CLK (.I(net384));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12201__CLK (.I(net384));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12344__CLK (.I(net385));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12169__CLK (.I(net385));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12207__CLK (.I(net385));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout384_I (.I(net385));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12178__CLK (.I(net386));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12175__CLK (.I(net386));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12173__CLK (.I(net386));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12172__CLK (.I(net386));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12171__CLK (.I(net386));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12177__CLK (.I(net387));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12176__CLK (.I(net387));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12168__CLK (.I(net387));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12179__CLK (.I(net387));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout386_I (.I(net387));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12180__CLK (.I(net388));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout387_I (.I(net388));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout385_I (.I(net388));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12184__CLK (.I(net389));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12183__CLK (.I(net389));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12182__CLK (.I(net389));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12181__CLK (.I(net389));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12167__CLK (.I(net389));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12188__CLK (.I(net390));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12185__CLK (.I(net390));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12165__CLK (.I(net390));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12164__CLK (.I(net390));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout389_I (.I(net391));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout390_I (.I(net391));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12260__CLK (.I(net391));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12166__CLK (.I(net391));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout391_I (.I(net392));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout388_I (.I(net392));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout392_I (.I(net393));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout382_I (.I(net393));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout393_I (.I(net394));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout367_I (.I(net394));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout394_I (.I(net395));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout338_I (.I(net395));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12196__CLK (.I(net396));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12197__CLK (.I(net396));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12143__CLK (.I(net396));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12141__CLK (.I(net396));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12140__CLK (.I(net396));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12152__CLK (.I(net398));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12144__CLK (.I(net398));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12199__CLK (.I(net398));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12195__CLK (.I(net398));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12139__CLK (.I(net398));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12200__CLK (.I(net399));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout398_I (.I(net399));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout397_I (.I(net399));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11998__CLK (.I(net400));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11997__CLK (.I(net400));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11996__CLK (.I(net400));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11517__CLK (.I(net400));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11516__CLK (.I(net400));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12151__CLK (.I(net401));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12090__CLK (.I(net401));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12089__CLK (.I(net401));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12000__CLK (.I(net401));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11999__CLK (.I(net401));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout400_I (.I(net402));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout401_I (.I(net402));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout399_I (.I(net402));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12091__CLK (.I(net403));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12194__CLK (.I(net403));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12193__CLK (.I(net403));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12138__CLK (.I(net403));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12137__CLK (.I(net403));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12126__CLK (.I(net405));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12098__CLK (.I(net405));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12130__CLK (.I(net405));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12128__CLK (.I(net405));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12121__CLK (.I(net405));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout405_I (.I(net406));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12125__CLK (.I(net406));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12124__CLK (.I(net406));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12123__CLK (.I(net406));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12122__CLK (.I(net406));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12127__CLK (.I(net407));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout406_I (.I(net407));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout403_I (.I(net407));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout404_I (.I(net407));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12005__CLK (.I(net408));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12004__CLK (.I(net408));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12096__CLK (.I(net408));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12095__CLK (.I(net408));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12094__CLK (.I(net408));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12129__CLK (.I(net410));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12097__CLK (.I(net410));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12081__CLK (.I(net410));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11983__CLK (.I(net410));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11981__CLK (.I(net410));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout410_I (.I(net412));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout411_I (.I(net412));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout408_I (.I(net412));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout409_I (.I(net412));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout412_I (.I(net413));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout407_I (.I(net413));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout413_I (.I(net414));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout402_I (.I(net414));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11701__CLK (.I(net415));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12003__CLK (.I(net415));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12002__CLK (.I(net415));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12001__CLK (.I(net415));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11718__CLK (.I(net415));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11726__CLK (.I(net416));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11710__CLK (.I(net416));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11709__CLK (.I(net416));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11702__CLK (.I(net416));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11717__CLK (.I(net417));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11712__CLK (.I(net417));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11696__CLK (.I(net417));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout415_I (.I(net417));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout416_I (.I(net417));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11862__CLK (.I(net420));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11858__CLK (.I(net420));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11857__CLK (.I(net420));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11427__CLK (.I(net420));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11840__CLK (.I(net421));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11846__CLK (.I(net421));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11844__CLK (.I(net421));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11839__CLK (.I(net421));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11704__CLK (.I(net421));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout421_I (.I(net423));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout422_I (.I(net423));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout419_I (.I(net423));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout420_I (.I(net423));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11708__CLK (.I(net425));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11700__CLK (.I(net425));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12011__CLK (.I(net425));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12010__CLK (.I(net425));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12009__CLK (.I(net425));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout428_I (.I(net429));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout425_I (.I(net429));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout426_I (.I(net429));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11522__CLK (.I(net430));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11521__CLK (.I(net430));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11525__CLK (.I(net430));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11520__CLK (.I(net430));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11519__CLK (.I(net430));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11845__CLK (.I(net432));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11843__CLK (.I(net432));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11842__CLK (.I(net432));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11526__CLK (.I(net432));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11524__CLK (.I(net432));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout431_I (.I(net433));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout432_I (.I(net433));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout429_I (.I(net433));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout433_I (.I(net434));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout424_I (.I(net434));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12135__CLK (.I(net436));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12133__CLK (.I(net436));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12132__CLK (.I(net436));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12131__CLK (.I(net436));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12082__CLK (.I(net436));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12136__CLK (.I(net438));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12134__CLK (.I(net438));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12088__CLK (.I(net438));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11985__CLK (.I(net438));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11984__CLK (.I(net438));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11955__CLK (.I(net440));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11954__CLK (.I(net440));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11953__CLK (.I(net440));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout438_I (.I(net440));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout439_I (.I(net440));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12104__CLK (.I(net441));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11957__CLK (.I(net441));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout440_I (.I(net442));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout441_I (.I(net442));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout436_I (.I(net442));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout437_I (.I(net442));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11947__CLK (.I(net444));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11946__CLK (.I(net444));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11945__CLK (.I(net444));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12102__CLK (.I(net444));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout443_I (.I(net444));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11973__CLK (.I(net446));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout445_I (.I(net446));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11969__CLK (.I(net446));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout446_I (.I(net447));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout444_I (.I(net447));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout447_I (.I(net448));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12099__CLK (.I(net448));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12083__CLK (.I(net448));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout448_I (.I(net449));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout442_I (.I(net449));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11722__CLK (.I(net450));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12018__CLK (.I(net450));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12017__CLK (.I(net450));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11714__CLK (.I(net450));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11713__CLK (.I(net450));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11721__CLK (.I(net452));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11698__CLK (.I(net452));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11697__CLK (.I(net452));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout450_I (.I(net452));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout451_I (.I(net452));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout453_I (.I(net455));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout454_I (.I(net455));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout452_I (.I(net455));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout456_I (.I(net457));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11918__CLK (.I(net457));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11911__CLK (.I(net457));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11910__CLK (.I(net457));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11903__CLK (.I(net457));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11894__CLK (.I(net458));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11886__CLK (.I(net458));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11917__CLK (.I(net458));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11912__CLK (.I(net458));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11904__CLK (.I(net458));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11902__CLK (.I(net459));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout458_I (.I(net459));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11896__CLK (.I(net459));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout457_I (.I(net459));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout459_I (.I(net460));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout455_I (.I(net460));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11908__CLK (.I(net461));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11949__CLK (.I(net461));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11948__CLK (.I(net461));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11944__CLK (.I(net461));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11943__CLK (.I(net461));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11941__CLK (.I(net462));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11940__CLK (.I(net462));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11936__CLK (.I(net462));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11909__CLK (.I(net462));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout465_I (.I(net467));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout466_I (.I(net467));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout461_I (.I(net467));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout462_I (.I(net467));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11900__CLK (.I(net468));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11893__CLK (.I(net468));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11892__CLK (.I(net468));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11885__CLK (.I(net468));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11884__CLK (.I(net468));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11899__CLK (.I(net471));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout470_I (.I(net471));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11906__CLK (.I(net471));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11905__CLK (.I(net471));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11898__CLK (.I(net471));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout471_I (.I(net472));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout469_I (.I(net472));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout472_I (.I(net473));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout467_I (.I(net473));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout473_I (.I(net474));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout460_I (.I(net474));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout475_I (.I(net476));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout435_I (.I(net476));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11860__CLK (.I(net477));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11859__CLK (.I(net477));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11822__CLK (.I(net477));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11816__CLK (.I(net477));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11815__CLK (.I(net477));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11838__CLK (.I(net478));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11833__CLK (.I(net478));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11832__CLK (.I(net478));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11831__CLK (.I(net478));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11817__CLK (.I(net478));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11767__CLK (.I(net479));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11760__CLK (.I(net479));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11759__CLK (.I(net479));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11752__CLK (.I(net479));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11751__CLK (.I(net479));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12021__CLK (.I(net481));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11769__CLK (.I(net481));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11768__CLK (.I(net481));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11761__CLK (.I(net481));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11753__CLK (.I(net481));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout481_I (.I(net483));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout482_I (.I(net483));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout479_I (.I(net483));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout480_I (.I(net483));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout483_I (.I(net484));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout477_I (.I(net484));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout478_I (.I(net484));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout485_I (.I(net487));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout486_I (.I(net487));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11837__CLK (.I(net487));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11836__CLK (.I(net487));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11530__CLK (.I(net488));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11529__CLK (.I(net488));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11527__CLK (.I(net488));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11534__CLK (.I(net488));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11533__CLK (.I(net488));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11531__CLK (.I(net489));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout488_I (.I(net489));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout487_I (.I(net489));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12026__CLK (.I(net490));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12025__CLK (.I(net490));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11770__CLK (.I(net490));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11762__CLK (.I(net490));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11754__CLK (.I(net490));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12262__CLK (.I(net491));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12261__CLK (.I(net491));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11771__CLK (.I(net491));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11763__CLK (.I(net491));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11755__CLK (.I(net491));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12307__CLK (.I(net492));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout491_I (.I(net492));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12027__CLK (.I(net492));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout490_I (.I(net492));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout492_I (.I(net493));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout489_I (.I(net493));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout493_I (.I(net494));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout484_I (.I(net494));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12023__CLK (.I(net495));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12292__CLK (.I(net495));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12291__CLK (.I(net495));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12046__CLK (.I(net495));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12045__CLK (.I(net495));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12162__CLK (.I(net497));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12189__CLK (.I(net497));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12187__CLK (.I(net497));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12186__CLK (.I(net497));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12161__CLK (.I(net497));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12192__CLK (.I(net498));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12191__CLK (.I(net498));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12190__CLK (.I(net498));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12163__CLK (.I(net498));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout497_I (.I(net499));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout498_I (.I(net499));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout495_I (.I(net499));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout496_I (.I(net499));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12289__CLK (.I(net500));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12407__CLK (.I(net500));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12304__CLK (.I(net500));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12303__CLK (.I(net500));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12047__CLK (.I(net500));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12332__CLK (.I(net501));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12331__CLK (.I(net501));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12290__CLK (.I(net501));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12305__CLK (.I(net502));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12287__CLK (.I(net502));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12286__CLK (.I(net502));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout500_I (.I(net502));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout501_I (.I(net502));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12284__CLK (.I(net504));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12283__CLK (.I(net504));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12330__CLK (.I(net504));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12329__CLK (.I(net504));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12328__CLK (.I(net504));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12285__CLK (.I(net505));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout504_I (.I(net505));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout502_I (.I(net505));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout503_I (.I(net505));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout505_I (.I(net506));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout499_I (.I(net506));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout506_I (.I(net507));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout494_I (.I(net507));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11847__CLK (.I(net508));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11764__CLK (.I(net508));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11851__CLK (.I(net508));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11850__CLK (.I(net508));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11849__CLK (.I(net508));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout509_I (.I(net510));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11878__CLK (.I(net510));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11854__CLK (.I(net510));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11853__CLK (.I(net510));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout510_I (.I(net511));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11872__CLK (.I(net511));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11871__CLK (.I(net511));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11528__CLK (.I(net511));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11774__CLK (.I(net512));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11766__CLK (.I(net512));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11758__CLK (.I(net512));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11757__CLK (.I(net512));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11756__CLK (.I(net512));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11773__CLK (.I(net514));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11772__CLK (.I(net514));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11765__CLK (.I(net514));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout512_I (.I(net514));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout513_I (.I(net514));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12265__CLK (.I(net515));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout514_I (.I(net515));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout511_I (.I(net515));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11863__CLK (.I(net516));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11877__CLK (.I(net516));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11876__CLK (.I(net516));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11870__CLK (.I(net516));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11869__CLK (.I(net516));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11867__CLK (.I(net519));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11865__CLK (.I(net519));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11875__CLK (.I(net519));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout518_I (.I(net519));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout519_I (.I(net520));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout516_I (.I(net520));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout517_I (.I(net520));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12268__CLK (.I(net521));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12267__CLK (.I(net521));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12266__CLK (.I(net521));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout520_I (.I(net521));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout521_I (.I(net522));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout515_I (.I(net522));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12309__CLK (.I(net523));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12335__CLK (.I(net523));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12334__CLK (.I(net523));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12308__CLK (.I(net523));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12288__CLK (.I(net523));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12317__CLK (.I(net524));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12310__CLK (.I(net524));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12279__CLK (.I(net525));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12327__CLK (.I(net525));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12326__CLK (.I(net525));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12282__CLK (.I(net525));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12281__CLK (.I(net525));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout525_I (.I(net527));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout526_I (.I(net527));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout523_I (.I(net527));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout524_I (.I(net527));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12271__CLK (.I(net530));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12270__CLK (.I(net530));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12269__CLK (.I(net530));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout528_I (.I(net530));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout529_I (.I(net530));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12322__CLK (.I(net532));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12321__CLK (.I(net532));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12320__CLK (.I(net532));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12319__CLK (.I(net532));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12278__CLK (.I(net532));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12277__CLK (.I(net533));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12276__CLK (.I(net533));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12275__CLK (.I(net533));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12274__CLK (.I(net533));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout532_I (.I(net534));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout533_I (.I(net534));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout530_I (.I(net534));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout531_I (.I(net534));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout534_I (.I(net535));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout527_I (.I(net535));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout535_I (.I(net536));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout522_I (.I(net536));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout536_I (.I(net537));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout507_I (.I(net537));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout537_I (.I(net538));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout476_I (.I(net538));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout538_I (.I(net539));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout395_I (.I(net539));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout539_I (.I(net540));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout269_I (.I(net540));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[18]_SE  (.I(net542));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[17]_SE  (.I(net542));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[16]_SE  (.I(net542));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[15]_SE  (.I(net542));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[14]_SE  (.I(net542));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[9]_SE  (.I(net544));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[13]_SE  (.I(net544));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[12]_SE  (.I(net544));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[11]_SE  (.I(net544));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[10]_SE  (.I(net544));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout544_I (.I(net546));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout545_I (.I(net546));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout542_I (.I(net546));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout543_I (.I(net546));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[31]_SE  (.I(net547));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[30]_SE  (.I(net547));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[28]_SE  (.I(net547));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[27]_SE  (.I(net547));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[3]_SE  (.I(net547));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[35]_SE  (.I(net549));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[34]_SE  (.I(net549));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[32]_SE  (.I(net549));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[8]_SE  (.I(net549));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout548_I (.I(net549));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout549_I (.I(net550));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[33]_SE  (.I(net550));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout547_I (.I(net550));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout550_I (.I(net551));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout546_I (.I(net551));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[40]_SE  (.I(net552));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[39]_SE  (.I(net552));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[38]_SE  (.I(net552));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[1]_SE  (.I(net552));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[0]_SE  (.I(net552));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[60]_SE  (.I(net554));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[67]_SE  (.I(net554));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[66]_SE  (.I(net554));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[65]_SE  (.I(net554));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[64]_SE  (.I(net554));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout554_I (.I(net556));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout555_I (.I(net556));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[63]_SE  (.I(net556));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[37]_SE  (.I(net556));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[36]_SE  (.I(net556));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout556_I (.I(net557));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout552_I (.I(net557));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout553_I (.I(net557));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[50]_SE  (.I(net558));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[49]_SE  (.I(net558));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[48]_SE  (.I(net558));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[47]_SE  (.I(net558));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[46]_SE  (.I(net558));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[69]_SE  (.I(net559));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[68]_SE  (.I(net559));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[45]_SE  (.I(net559));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[44]_SE  (.I(net559));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[43]_SE  (.I(net559));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[56]_SE  (.I(net561));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[55]_SE  (.I(net561));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[54]_SE  (.I(net561));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[53]_SE  (.I(net561));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[52]_SE  (.I(net561));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[58]_SE  (.I(net562));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout561_I (.I(net562));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[59]_SE  (.I(net562));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[57]_SE  (.I(net562));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout562_I (.I(net563));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout559_I (.I(net563));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout560_I (.I(net563));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout563_I (.I(net564));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout557_I (.I(net564));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout564_I (.I(net565));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout551_I (.I(net565));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1758 ();
 assign io_oeb[0] = net566;
 assign io_oeb[1] = net567;
 assign io_oeb[2] = net568;
 assign io_oeb[3] = net569;
 assign io_oeb[4] = net570;
 assign io_out[2] = net571;
 assign io_out[3] = net572;
 assign io_out[4] = net573;
endmodule

