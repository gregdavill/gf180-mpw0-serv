* NGSPICE file created from serv_0.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__sdffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__sdffq_1 D SE SI CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyd_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyd_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_4 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnq_1 D CLKN Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_12 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_ip_sram__sram256x8m8wm1 abstract view
.subckt gf180mcu_fd_ip_sram__sram256x8m8wm1 A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7]
+ CEN CLK D[0] D[1] D[2] D[3] D[4] D[5] D[6] D[7] GWEN Q[0] Q[1] Q[2] Q[3] Q[4] Q[5]
+ Q[6] Q[7] WEN[0] WEN[1] WEN[2] WEN[3] WEN[4] WEN[5] WEN[6] WEN[7] VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_2 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_3 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

.subckt serv_0 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_oeb[0] io_oeb[1] io_oeb[2]
+ io_oeb[3] io_oeb[4] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] vdd vss
XFILLER_41_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3155_ _0013_ net65 u_cpu.cpu.alu.add_cy_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout56_I net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3086_ _0111_ net68 u_cpu.cpu.genblk3.csr.timer_irq_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2106_ u_cpu.cpu.state.init_done _0287_ _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2037_ _1045_ u_cpu.cpu.state.stage_two_req _0254_ _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_63_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[45\]_SE net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2939_ _0985_ _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2182__A2 _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3132__CLK net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1693__A1 _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2245__I0 u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[34\] u_arbiter.i_wb_cpu_rdt\[31\] net144 u_arbiter.i_wb_cpu_dbus_dat\[28\]
+ net30 u_scanchain_local.module_data_in\[34\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_64_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[68\]_SE net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3005__CLK net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2724_ _0845_ _0124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2655_ u_cpu.cpu.immdec.imm19_12_20\[6\] _0568_ _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1606_ _1080_ _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3155__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2586_ _0732_ _0731_ _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout116 net122 net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout127 net128 net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout105 net109 net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout138 net139 net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout149 net150 net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_80_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3207_ _0211_ net52 u_cpu.rf_ram_if.rdata1\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3138_ _0160_ net112 u_cpu.cpu.ctrl.o_ibus_adr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1675__A1 _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3069_ _0094_ net61 u_cpu.cpu.immdec.imm30_25\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1978__A2 _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1666__A1 _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3028__CLK net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout106_I net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2440_ _0598_ _0599_ _0536_ _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_142_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2371_ _0513_ _0509_ _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2082__A1 _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout19_I net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2707_ u_arbiter.i_wb_cpu_dbus_adr\[6\] u_arbiter.i_wb_cpu_dbus_adr\[7\] _0831_ _0836_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2385__A2 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2137__A2 _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2638_ _0542_ _0778_ _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2569_ _0415_ _0485_ _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2860__A3 _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2073__A1 _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1958__S _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1820__A1 _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2923__I1 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1887__A1 _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2687__I0 u_arbiter.i_wb_cpu_rdt\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1940_ _1353_ _0021_ _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1667__I _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1811__A1 _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1871_ _1293_ _1282_ _1295_ _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_35_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2699__S _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2119__A2 _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2423_ _0442_ _0582_ _0583_ _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2354_ _1079_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[11\] _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_9_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2285_ u_arbiter.i_wb_cpu_rdt\[1\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\] _1079_
+ _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1869__A1 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2530__A2 _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2818__B1 _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1688__S _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2046__A1 u_arbiter.i_wb_cpu_dbus_dat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2597__A2 _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3216__CLK net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2070_ _0246_ _0280_ _0281_ _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_75_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2972_ u_cpu.cpu.ctrl.i_iscomp _0413_ _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2037__A1 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2588__A2 _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1923_ u_cpu.rf_ram_if.wdata0_r\[6\] u_cpu.rf_ram_if.wdata1_r\[6\] _1341_ _1349_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1854_ _1282_ _1295_ _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1785_ _1208_ _1227_ _1228_ _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2760__A2 _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2021__I _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2406_ _0254_ _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_fanout86_I net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2337_ _0426_ _0433_ _0501_ _0503_ _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2268_ _0423_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\] _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1866__A4 _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2199_ u_arbiter.i_wb_cpu_dbus_dat\[19\] _0375_ _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2579__A2 _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2200__A1 u_arbiter.i_wb_cpu_rdt\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2503__A2 _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2267__A1 _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2019__A1 u_cpu.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xu_scanchain_local.scan_flop\[64\] u_scanchain_local.module_data_in\[63\] net148 u_arbiter.o_wb_cpu_adr\[26\]
+ net34 u_scanchain_local.module_data_in\[64\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XPHY_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1570_ _1048_ _1031_ _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_4_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3171_ _0192_ net91 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2776__I _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2122_ _0322_ _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2053_ _0255_ _0269_ _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2955_ u_cpu.cpu.genblk3.csr.mcause31 _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_124_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1906_ _1339_ _0023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2886_ _0932_ _0949_ _0950_ _0952_ _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1837_ _1275_ _1278_ _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1768_ u_cpu.rf_ram_if.rcnt\[0\] _1021_ _1022_ u_cpu.rf_ram_if.wen0_r _1212_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_132_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1699_ _1155_ _1156_ _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3061__CLK net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2972__A2 _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput7 net7 io_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_114_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2529__C _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2740_ u_arbiter.i_wb_cpu_dbus_adr\[21\] u_arbiter.i_wb_cpu_dbus_adr\[22\] _0849_
+ _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_fanout136_I net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2671_ _0415_ _0774_ _0807_ _0808_ _0799_ _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__2963__A2 _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1622_ u_arbiter.i_wb_cpu_dbus_adr\[3\] _1091_ _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1553_ _1031_ _1032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_141_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2479__A1 _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3154_ _0176_ net81 u_cpu.cpu.ctrl.o_ibus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3085_ _0110_ net75 u_cpu.cpu.immdec.imm31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2105_ _0307_ _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2036_ _0253_ _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_fanout49_I net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3084__CLK net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2938_ u_arbiter.i_wb_cpu_rdt\[31\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\]
+ _0252_ _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2403__A1 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2869_ _0799_ _0936_ _0561_ _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2167__B1 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2890__A1 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[27\] u_arbiter.i_wb_cpu_rdt\[24\] net130 u_arbiter.i_wb_cpu_dbus_dat\[21\]
+ net16 u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_69_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1684__A2 _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2881__A1 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2633__A1 _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2723_ u_arbiter.i_wb_cpu_dbus_adr\[13\] u_arbiter.i_wb_cpu_dbus_adr\[14\] _0843_
+ _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2654_ _0474_ _0782_ _0793_ _0477_ _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1605_ _1079_ _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2585_ u_cpu.cpu.immdec.imm31 _1222_ _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xfanout117 net121 net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
Xfanout128 net129 net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout106 net109 net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout139 net140 net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[12\]_SE net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3206_ u_cpu.rf_ram_if.wtrig0 net51 u_cpu.rf_ram_if.genblk1.wtrig0_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3137_ _0159_ net112 u_cpu.cpu.ctrl.o_ibus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2872__A1 _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3068_ _0093_ net60 u_cpu.cpu.immdec.imm24_20\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2019_ u_cpu.cpu.immdec.imm11_7\[1\] u_cpu.cpu.immdec.imm11_7\[2\] u_cpu.cpu.immdec.imm11_7\[3\]
+ u_cpu.cpu.immdec.imm11_7\[0\] _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_24_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1978__A3 _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[23\]_CLK net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[38\]_CLK net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[35\]_SE net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2370_ _0468_ _0534_ _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2606__A1 _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2606__B2 _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2082__A2 _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3122__CLK net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2706_ _0835_ _0116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2637_ _0528_ _0508_ _0768_ _0777_ _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_12_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2568_ _0457_ _0715_ _0583_ _0578_ _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2499_ _0546_ _0650_ _0652_ _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1648__A2 _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2627__C _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2073__A2 _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1820__A2 _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1773__I u_cpu.cpu.bufreg2.i_cnt_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2687__I1 u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3145__CLK net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1811__A2 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1870_ _1301_ _1306_ _1309_ _1311_ _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_35_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2221__C1 _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2779__I _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1575__A1 _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2422_ _0471_ _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2353_ _0518_ _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2284_ _0430_ u_arbiter.i_wb_cpu_rdt\[0\] _0452_ _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_42_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout31_I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2212__C1 _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1999_ _1264_ _0224_ _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1593__I _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3018__CLK net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2530__A3 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[1\]_CLK net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_93_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2046__A2 _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2373__B _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2971_ _1006_ _1007_ _1008_ _1009_ _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_124_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1922_ _1348_ u_cpu.rf_ram.i_wdata\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1853_ _1287_ _1294_ _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1784_ _1207_ u_cpu.cpu.alu.add_cy_r _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout8 net10 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_131_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2405_ _0215_ _0515_ _0567_ _0083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1720__A1 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2336_ _0470_ _0502_ _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout79_I net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2267_ _0430_ u_arbiter.i_wb_cpu_rdt\[6\] _0435_ _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_66_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2198_ _0379_ _0381_ _0062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1789__S _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2200__A2 _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2267__A2 u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_scanchain_local.scan_flop\[57\] u_scanchain_local.module_data_in\[56\] net142 u_arbiter.o_wb_cpu_adr\[19\]
+ net28 u_scanchain_local.module_data_in\[57\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__2550__C _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2122__I _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3170_ _0191_ net90 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1702__A1 _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2121_ _0320_ _0313_ _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2052_ u_cpu.cpu.state.init_done _1046_ _0218_ _0268_ _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_63_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2954_ _0993_ _0989_ _0996_ _1261_ _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2885_ _0542_ _0703_ _0951_ _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1905_ u_cpu.rf_ram.rdata\[6\] u_cpu.rf_ram.data\[6\] _1203_ _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1836_ u_cpu.cpu.state.stage_two_req _1277_ _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1767_ _1200_ _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_117_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1698_ u_cpu.cpu.ctrl.o_ibus_adr\[18\] u_cpu.cpu.ctrl.o_ibus_adr\[17\] u_cpu.cpu.ctrl.o_ibus_adr\[16\]
+ _1145_ _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_44_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2497__A2 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2319_ _0486_ _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3206__CLK net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2732__I0 u_arbiter.i_wb_cpu_dbus_adr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[2\] net12 net135 u_arbiter.i_wb_cpu_dbus_sel\[0\] net22
+ u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_37_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2670_ _0524_ _0741_ _0554_ _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2963__A3 _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1621_ u_cpu.cpu.ctrl.o_ibus_adr\[3\] _1086_ _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_67_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1552_ u_cpu.cpu.branch_op _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_67_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3153_ _0175_ net108 u_cpu.cpu.ctrl.o_ibus_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2479__A2 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input3_I io_in[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2104_ _1246_ _1290_ _0039_ _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_36_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3084_ _0109_ net60 u_cpu.cpu.immdec.imm19_12_20\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2035_ _0251_ u_arbiter.i_wb_cpu_ibus_adr\[1\] _0252_ _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2651__A2 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2937_ _0984_ _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout8_I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2868_ _0462_ _0741_ _0786_ _0935_ _0554_ _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_136_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2799_ _0891_ _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2167__A1 u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2167__B2 u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1819_ _1052_ _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2697__I _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2714__I0 u_arbiter.i_wb_cpu_dbus_adr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[9\]_SE net136 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2365__C _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2330__A1 _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1841__B1 _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2722_ _0844_ _0123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2653_ _0783_ _0784_ _0496_ _0792_ _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1604_ _1078_ _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2584_ _1320_ _0297_ _0222_ _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xfanout118 net121 net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout129 net133 net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout107 net108 net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_86_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3051__CLK net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3205_ u_cpu.cpu.o_wdata0 net47 u_cpu.rf_ram_if.wdata0_r\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3136_ _0158_ net111 u_cpu.cpu.ctrl.o_ibus_adr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout61_I net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3067_ _0092_ net47 u_cpu.cpu.immdec.imm24_20\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2018_ _1053_ _0219_ u_cpu.cpu.o_wen1 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_24_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2560__B2 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1666__A3 _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3074__CLK net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2303__A1 _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1901__I1 u_cpu.rf_ram.data\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2705_ u_arbiter.i_wb_cpu_dbus_adr\[5\] u_arbiter.i_wb_cpu_dbus_adr\[6\] _0831_ _0835_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2636_ _0769_ _0743_ _0776_ _0622_ _0496_ _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__2917__I0 u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2567_ _0251_ u_arbiter.i_wb_cpu_rdt\[13\] _0714_ _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2542__A1 _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2498_ _0526_ _0651_ _0607_ _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_59_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3119_ _0143_ net77 u_cpu.cpu.bufreg.lsb\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3097__CLK net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1584__A2 _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2908__I0 u_arbiter.i_wb_cpu_rdt\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3193__D _0021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2533__A1 _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2221__B1 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2221__C2 u_arbiter.i_wb_cpu_dbus_dat\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout111_I net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2524__A1 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2421_ _0494_ _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2352_ _0448_ _0459_ _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2283_ _0427_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\] _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[22\]_CLK net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_u_scanchain_local.scan_flop\[37\]_CLK net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout24_I net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2212__B1 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1998_ _1271_ _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2619_ u_cpu.cpu.immdec.imm19_12_20\[3\] _0505_ _0757_ _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_47_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2515__A1 _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2818__A2 _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_93_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_93_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[25\]_SE net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2203__B1 _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[32\]_SI u_arbiter.i_wb_cpu_dbus_dat\[26\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3112__CLK net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2970_ u_cpu.cpu.genblk3.csr.mstatus_mie _1000_ _1007_ _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1895__S _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1921_ u_cpu.rf_ram_if.wdata0_r\[5\] u_cpu.rf_ram_if.wdata1_r\[5\] _1341_ _1348_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1852_ _1289_ _1291_ _1293_ _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1783_ _1206_ _1226_ _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xfanout9 net10 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_118_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2404_ _0467_ _0561_ _0566_ _0514_ _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2335_ _0480_ _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2266_ _0423_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[6\] _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_66_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2197_ u_arbiter.i_wb_cpu_rdt\[17\] _0380_ _0371_ u_arbiter.i_wb_cpu_dbus_dat\[17\]
+ _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_u_scanchain_local.scan_flop\[48\]_SE net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3135__CLK net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2019__A3 u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1778__A2 _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2975__A1 _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1702__A2 _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2120_ _0320_ _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2051_ _1310_ _0265_ _0267_ _1033_ _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_63_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2953_ _1039_ _1050_ _0989_ _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3008__CLK net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1904_ _1338_ _0022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2884_ _0608_ _0449_ _0509_ _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1835_ _1028_ u_arbiter.i_wb_cpu_dbus_dat\[5\] _1276_ u_cpu.cpu.state.init_done _1277_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__3158__CLK net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[0\]_CLK net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1766_ u_cpu.rf_ram.data\[0\] _1200_ _1201_ _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_1697_ u_cpu.cpu.ctrl.o_ibus_adr\[19\] _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_fanout91_I net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2318_ _0440_ _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_44_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2249_ u_arbiter.i_wb_cpu_rdt\[7\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[7\] _0416_
+ _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_54_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2957__A1 _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2223__I u_arbiter.i_wb_cpu_dbus_dat\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2248__I0 u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2963__A4 _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1620_ _1093_ _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2176__A2 _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1551_ u_cpu.cpu.decode.opcode\[2\] _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_28_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3221_ u_cpu.cpu.o_wen1 net55 u_cpu.rf_ram_if.wen1_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2723__I1 u_arbiter.i_wb_cpu_dbus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3152_ _0174_ net117 u_cpu.cpu.ctrl.o_ibus_adr\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2103_ _0296_ _0306_ _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3083_ _0108_ net48 u_cpu.cpu.immdec.imm19_12_20\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2034_ net12 _1073_ _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__2636__B1 _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2308__I _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2936_ u_arbiter.i_wb_cpu_rdt\[30\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[14\]
+ _0979_ _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1611__A1 _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2867_ _0421_ _0631_ _0582_ _0486_ _0741_ _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_11_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1818_ _1234_ _1260_ _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2798_ u_cpu.cpu.ctrl.o_ibus_adr\[8\] _0885_ _0887_ u_cpu.cpu.ctrl.o_ibus_adr\[9\]
+ _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2167__A2 _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1749_ _1074_ _1195_ _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2330__A2 _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1967__I _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1841__B2 _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout141_I net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2721_ u_arbiter.i_wb_cpu_dbus_adr\[12\] u_arbiter.i_wb_cpu_dbus_adr\[13\] _0843_
+ _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2652_ _0788_ _0791_ _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1603_ u_cpu.cpu.genblk1.align.ctrl_misal _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2583_ u_cpu.cpu.immdec.imm19_12_20\[0\] _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout119 net121 net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout108 net109 net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_3204_ u_cpu.rf_ram_if.wdata0_r\[6\] net47 u_cpu.rf_ram_if.wdata0_r\[5\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3135_ _0157_ net111 u_cpu.cpu.ctrl.o_ibus_adr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout54_I net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3066_ _0091_ net49 u_cpu.cpu.immdec.imm24_20\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2017_ _0239_ _0240_ _0238_ _0015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2919_ u_arbiter.i_wb_cpu_rdt\[22\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[6\]
+ _0973_ _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2699__I0 u_arbiter.i_wb_cpu_dbus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2076__A1 _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3219__CLK net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[32\] u_arbiter.i_wb_cpu_rdt\[29\] net144 u_arbiter.i_wb_cpu_dbus_dat\[26\]
+ net30 u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__2000__A1 _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2303__A2 _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1814__A1 _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2704_ _0834_ _0115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2635_ _0775_ _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2917__I1 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2566_ _0589_ u_arbiter.i_wb_cpu_rdt\[29\] _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__2542__A2 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2497_ _0425_ _0543_ _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3118_ _0014_ net74 u_cpu.cpu.bufreg.c_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3049_ _0074_ net102 u_arbiter.i_wb_cpu_dbus_dat\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2058__A1 u_cpu.raddr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1805__A1 u_cpu.cpu.decode.op26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2908__I1 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1895__I1 u_cpu.rf_ram.data\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2049__A1 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2406__I _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3041__CLK net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout90 net96 net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_35_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2221__A1 u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2141__I _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout104_I net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2420_ _0426_ _0449_ _0580_ _0442_ _0433_ _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__1980__B1 _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3191__CLK net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2351_ _0516_ _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2282_ _0426_ _0450_ _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_81_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2316__I _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout17_I net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1997_ _1264_ _0222_ _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2212__A1 u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2618_ u_cpu.cpu.immdec.imm19_12_20\[2\] _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_115_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2549_ _0487_ _0631_ _0433_ _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2654__C _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3064__CLK net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2670__B _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2203__A1 u_arbiter.i_wb_cpu_rdt\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1876__S0 u_cpu.cpu.bufreg.lsb\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1920_ _1347_ u_cpu.rf_ram.i_wdata\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1851_ _1264_ _1292_ _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1782_ _1209_ _1215_ _1216_ _1225_ _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2403_ _0517_ _0565_ _0503_ _0561_ _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2334_ _0500_ _0444_ _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_130_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2265_ _0429_ _0433_ _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_93_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2196_ _0338_ _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_77_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3087__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2681__A1 _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2681__B2 _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2474__C _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2433__A1 _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2197__B1 _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2710__S _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1711__A3 _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2672__A1 _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2019__A4 u_cpu.cpu.immdec.imm11_7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2424__A1 _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1795__I _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[21\]_CLK net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[36\]_CLK net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2050_ _0266_ _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2663__A1 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2952_ _0992_ _0989_ _0995_ _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_37_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1903_ u_cpu.rf_ram.rdata\[5\] u_cpu.rf_ram.data\[5\] _1333_ _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2883_ u_cpu.cpu.immdec.imm11_7\[2\] _0932_ _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1834_ _1035_ _1030_ _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA_u_scanchain_local.scan_flop\[20\]_D u_arbiter.i_wb_cpu_rdt\[17\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1765_ u_arbiter.i_wb_cpu_dbus_we _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_1696_ _1154_ u_arbiter.o_wb_cpu_adr\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[15\]_SE net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout84_I net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2317_ _0484_ _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2248_ u_arbiter.i_wb_cpu_rdt\[9\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[9\] _0416_
+ _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2179_ _0320_ _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2654__A1 _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2705__S _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[22\]_SI u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3102__CLK net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[11\]_D u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2893__A1 _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2645__A1 _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[62\] u_scanchain_local.module_data_in\[61\] net145 u_arbiter.o_wb_cpu_adr\[24\]
+ net33 u_scanchain_local.module_data_in\[62\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA_u_scanchain_local.scan_flop\[9\]_D u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1550_ _1028_ _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_119_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[38\]_SE net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3220_ u_cpu.cpu.o_wen0 net55 u_cpu.rf_ram_if.wen0_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3151_ _0173_ net118 u_cpu.cpu.ctrl.o_ibus_adr\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1687__A2 _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2102_ _0297_ _0305_ _0032_ _1266_ _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__2884__A1 _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3082_ _0107_ net48 u_cpu.cpu.immdec.imm19_12_20\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2033_ _0250_ _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2636__B2 _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2935_ _0983_ _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2866_ _0695_ _0434_ _0501_ _0534_ _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__2324__I _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1817_ _1235_ _1242_ _1257_ _1259_ _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_2797_ _0890_ _0152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1748_ u_cpu.cpu.ctrl.o_ibus_adr\[30\] u_cpu.cpu.ctrl.o_ibus_adr\[29\] _1191_ _1195_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_144_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1679_ _1140_ _1137_ _1141_ _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2875__B2 _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2875__A1 _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2627__A1 _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1850__A2 _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1669__A2 _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2866__A1 _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3148__CLK net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2720_ _1288_ _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_fanout134_I net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2651_ _0656_ _0503_ _0790_ _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_34_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1602_ _1077_ u_arbiter.o_wb_cpu_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2582_ u_cpu.cpu.immdec.imm30_25\[5\] _0688_ _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout109 net110 net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_10_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3203_ u_cpu.rf_ram_if.wdata0_r\[5\] net44 u_cpu.rf_ram_if.wdata0_r\[4\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3134_ _0156_ net111 u_cpu.cpu.ctrl.o_ibus_adr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2319__I _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2609__A1 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3065_ _0090_ net57 u_cpu.cpu.immdec.imm24_20\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2016_ _1325_ _1326_ _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2255__S _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout47_I net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2763__B _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1832__A2 _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2918_ _0974_ _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1596__A1 _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2849_ _0920_ _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_12_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2784__B1 _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1587__A1 _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[25\] u_arbiter.i_wb_cpu_rdt\[22\] net129 u_arbiter.i_wb_cpu_dbus_dat\[19\]
+ net15 u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_29_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2311__I0 u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1814__A2 _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2703_ u_arbiter.i_wb_cpu_dbus_adr\[4\] u_arbiter.i_wb_cpu_dbus_adr\[5\] _0831_ _0834_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2634_ _0771_ _0772_ _0774_ _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_12_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2565_ _0710_ _0712_ _0713_ _0097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_12_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1750__A1 u_arbiter.i_wb_cpu_dbus_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2496_ _0608_ _0607_ _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3117_ _0142_ net81 u_arbiter.i_wb_cpu_dbus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3048_ _0073_ net102 u_arbiter.i_wb_cpu_dbus_dat\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2493__B _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1584__A4 _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2518__B1 _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2387__C _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2049__A2 _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout91 net95 net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_35_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout80 net83 net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_70_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2221__A2 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1980__B2 _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2350_ _0429_ _0432_ _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2281_ _0434_ _0449_ _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1799__A1 _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1996_ u_cpu.cpu.decode.opcode\[1\] _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2212__A2 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2617_ _0759_ _0756_ _0760_ _0560_ _0102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_138_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2548_ _0420_ _0494_ _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2479_ _0588_ _0616_ _0633_ _0636_ _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_29_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3209__CLK net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_58_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_93_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2203__A2 _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2242__I _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1714__A1 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1876__S1 _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2442__A2 _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1850_ _1048_ _1271_ _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1781_ _1204_ _1224_ _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_129_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1991__I _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2402_ _0486_ _0543_ _0519_ _0563_ _0564_ _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_130_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2753__I0 u_arbiter.i_wb_cpu_dbus_adr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2333_ _0493_ _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2264_ _0432_ _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2195_ u_arbiter.i_wb_cpu_dbus_dat\[18\] _0375_ _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2528__S _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2130__A1 u_arbiter.i_wb_cpu_rdt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2681__A2 _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2433__A2 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2490__C _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2197__A1 u_arbiter.i_wb_cpu_rdt\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2197__B2 u_arbiter.i_wb_cpu_dbus_dat\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1979_ u_cpu.cpu.immdec.imm11_7\[2\] _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3031__CLK net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2672__A2 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_45_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3181__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2424__A2 _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2415__A2 _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2951_ _1047_ _1033_ _0988_ _0994_ _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_76_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1902_ _1337_ _0021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2882_ u_cpu.cpu.immdec.imm11_7\[3\] _0638_ _0498_ _0948_ _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1833_ _1269_ _1274_ _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1764_ _1207_ u_cpu.cpu.alu.add_cy_r _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1695_ u_arbiter.i_wb_cpu_dbus_adr\[18\] _1153_ _1074_ _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2610__I _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3054__CLK net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2316_ _0483_ _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2766__B _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout77_I net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2247_ _0248_ _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2178_ _0366_ _0367_ _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2654__A2 _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2342__A1 _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xu_scanchain_local.scan_flop\[55\] u_scanchain_local.module_data_in\[54\] net143 u_arbiter.o_wb_cpu_adr\[17\]
+ net29 u_scanchain_local.module_data_in\[55\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2430__I _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2581__B2 _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2581__A1 _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3150_ _0172_ net118 u_cpu.cpu.ctrl.o_ibus_adr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2884__A2 _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2101_ _1235_ _0304_ _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3081_ _0106_ net47 u_cpu.cpu.immdec.imm19_12_20\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2032_ _0249_ _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_36_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2934_ u_arbiter.i_wb_cpu_rdt\[29\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[13\]
+ _0979_ _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2865_ _1218_ _0932_ _0933_ _0749_ _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1816_ _1258_ _1235_ _1241_ _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2796_ u_cpu.cpu.ctrl.o_ibus_adr\[7\] _0885_ _0887_ u_cpu.cpu.ctrl.o_ibus_adr\[8\]
+ _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1747_ u_cpu.cpu.ctrl.o_ibus_adr\[29\] _1191_ u_cpu.cpu.ctrl.o_ibus_adr\[30\] _1194_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_11_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1678_ _1140_ _1137_ _1093_ _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2875__A2 _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[20\]_CLK net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2627__A2 _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2716__S _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[35\]_CLK net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2938__I0 u_arbiter.i_wb_cpu_rdt\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2866__A2 _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_scanchain_local.scan_flop\[0\] net3 net139 u_arbiter.o_wb_cpu_cyc net25 u_cpu.cpu.genblk3.csr.i_mtip
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_92_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_fanout127_I net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2650_ _0421_ _0434_ _0789_ _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_34_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1601_ u_arbiter.i_wb_cpu_ibus_adr\[1\] _1073_ _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2581_ _0510_ _0723_ _0727_ _0514_ _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_45_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3202_ u_cpu.rf_ram_if.wdata0_r\[4\] net41 u_cpu.rf_ram_if.wdata0_r\[3\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input1_I io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2857__A2 _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3133_ _0155_ net113 u_cpu.cpu.ctrl.o_ibus_adr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_u_scanchain_local.scan_flop\[12\]_SI u_arbiter.i_wb_cpu_dbus_dat\[6\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3064_ _0089_ net57 u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2015_ _1071_ u_cpu.cpu.ctrl.pc_plus_4_cy_r _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2917_ u_arbiter.i_wb_cpu_rdt\[21\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\]
+ _0973_ _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2848_ u_cpu.cpu.ctrl.o_ibus_adr\[29\] _0876_ _0915_ u_cpu.cpu.ctrl.o_ibus_adr\[30\]
+ _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2779_ _0879_ _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2848__A2 _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2673__C _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[28\]_SE net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1587__A2 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2536__A1 _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3115__CLK net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[18\] u_arbiter.i_wb_cpu_rdt\[15\] net127 u_arbiter.i_wb_cpu_dbus_dat\[12\]
+ net13 u_arbiter.i_wb_cpu_rdt\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_2_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2472__B1 _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2155__I _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2702_ _0833_ _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2633_ _0444_ _0773_ _0608_ _0480_ _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2564_ _0477_ _0561_ _0707_ _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_12_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2527__A1 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1750__A2 _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2495_ u_arbiter.i_wb_cpu_rdt\[23\] u_arbiter.i_wb_cpu_rdt\[7\] _1081_ _0649_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3116_ _0141_ net82 u_arbiter.i_wb_cpu_dbus_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2774__B net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3047_ _0072_ net102 u_arbiter.i_wb_cpu_dbus_dat\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2215__B1 _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2518__B2 _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1741__A2 _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2206__B1 _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout92 net95 net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout81 net83 net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout70 net71 net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_35_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2509__A1 _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2578__C _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2280_ _0444_ _0448_ _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_81_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1995_ _1209_ _1075_ u_arbiter.o_wb_cpu_we vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_140_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2616_ u_cpu.cpu.immdec.imm19_12_20\[2\] _0505_ _0757_ _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2547_ _0695_ _0557_ _0696_ _0664_ _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2478_ _0598_ _0635_ _0537_ _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_93_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2987__A1 _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2523__I _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2679__B _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2278__I0 u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1780_ _1217_ _1220_ _1221_ _1223_ _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_115_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2401_ _0552_ _0483_ _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1705__A2 _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2902__A1 u_arbiter.i_wb_cpu_ack vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2332_ _0491_ _0495_ _0498_ _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2263_ _0430_ u_arbiter.i_wb_cpu_rdt\[1\] _0431_ _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_46_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2194_ _0378_ _0061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2130__A2 _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout22_I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1641__A1 _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2197__A2 _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1978_ _1350_ _1066_ _1202_ _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_101_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2121__A2 _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2409__B1 _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1632__A1 _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_61_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2428__I _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2950_ _0993_ _1262_ _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2820__B1 _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1623__A1 _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2881_ _0603_ _0944_ _0947_ _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1901_ u_cpu.rf_ram.rdata\[4\] u_cpu.rf_ram.data\[4\] _1333_ _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1832_ _1230_ _1273_ _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1763_ u_cpu.cpu.alu.i_rs1 _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1694_ u_cpu.cpu.ctrl.o_ibus_adr\[18\] _1151_ _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_125_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2315_ _0480_ _0482_ _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2766__C _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2246_ u_arbiter.i_wb_cpu_rdt\[10\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[10\]
+ _0248_ _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2177_ u_arbiter.i_wb_cpu_rdt\[11\] _0364_ _0348_ u_arbiter.i_wb_cpu_dbus_dat\[11\]
+ _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[61\]_SE net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2590__A2 _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2022__B _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2912__S _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xu_scanchain_local.scan_flop\[48\] u_scanchain_local.module_data_in\[47\] net141 u_arbiter.o_wb_cpu_adr\[10\]
+ net27 u_scanchain_local.module_data_in\[48\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_67_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2581__A2 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1771__B u_cpu.rf_ram.regzero vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2100_ _0298_ _0302_ _0303_ _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3080_ _0105_ net57 u_cpu.cpu.csr_imm vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2031_ _0248_ _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_130_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2933_ _0982_ _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2864_ u_cpu.cpu.immdec.imm11_7\[1\] _0638_ _0932_ _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2795_ _0889_ _0151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1815_ _1035_ _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1746_ _1111_ _1192_ _1193_ u_arbiter.o_wb_cpu_adr\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3021__CLK net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1677_ u_cpu.cpu.ctrl.o_ibus_adr\[14\] _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3171__CLK net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2229_ u_arbiter.i_wb_cpu_rdt\[28\] _0338_ _0390_ u_arbiter.i_wb_cpu_dbus_dat\[28\]
+ _0346_ u_arbiter.i_wb_cpu_dbus_dat\[29\] _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_2_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1901__S _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1835__A1 _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2732__S _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2315__A2 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2866__A3 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2079__A1 _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1826__A1 u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2642__S _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1600_ _1076_ u_arbiter.o_wb_cpu_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2580_ _0620_ _0726_ _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3194__CLK net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3201_ u_cpu.rf_ram_if.wdata0_r\[3\] net40 u_cpu.rf_ram_if.wdata0_r\[2\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3132_ _0154_ net103 u_cpu.cpu.ctrl.o_ibus_adr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3063_ _0088_ net75 u_cpu.cpu.decode.op26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2014_ _0234_ _0236_ _0238_ _0016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1817__A1 _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2916_ _0252_ _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2847_ _0919_ _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2778_ _0878_ _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1729_ _1174_ _1179_ _1180_ u_arbiter.o_wb_cpu_adr\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1808__A1 _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2233__A1 u_arbiter.i_wb_cpu_rdt\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2000__A4 _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1605__I _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2472__A1 _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2472__B2 _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2701_ u_arbiter.i_wb_cpu_dbus_adr\[3\] u_arbiter.i_wb_cpu_dbus_adr\[4\] _0831_ _0833_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2632_ _0424_ _0493_ _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2563_ u_cpu.cpu.immdec.imm30_25\[3\] _0685_ _0711_ u_cpu.cpu.immdec.imm30_25\[4\]
+ _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__2527__A2 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2494_ _0647_ _0642_ _0648_ _0614_ _0091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_96_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[34\]_CLK net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3115_ _0140_ net108 u_arbiter.i_wb_cpu_dbus_adr\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3046_ _0071_ net102 u_arbiter.i_wb_cpu_dbus_dat\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout52_I net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[49\]_CLK net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2215__A1 u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2766__A2 _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2965__B _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2256__I _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2454__A1 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2206__A1 u_arbiter.i_wb_cpu_rdt\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout82 net83 net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_35_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout71 net72 net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_23_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout60 net62 net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
Xfanout93 net95 net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_11_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2509__A2 _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_scanchain_local.scan_flop\[30\] u_arbiter.i_wb_cpu_rdt\[27\] net131 u_arbiter.i_wb_cpu_dbus_dat\[24\]
+ net17 u_arbiter.i_wb_cpu_rdt\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_81_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3202__D u_cpu.rf_ram_if.wdata0_r\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1994_ _0217_ _0221_ _1094_ u_arbiter.o_wb_cpu_cyc vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2615_ u_cpu.cpu.immdec.imm19_12_20\[1\] _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_86_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[18\]_SE net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2546_ u_arbiter.i_wb_cpu_rdt\[27\] u_arbiter.i_wb_cpu_rdt\[11\] _1082_ _0696_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_47_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2477_ _0466_ _0546_ _0448_ _0616_ _0634_ _0622_ _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_96_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2684__A1 _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3029_ _0054_ net94 u_arbiter.i_wb_cpu_dbus_dat\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2436__A1 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3105__CLK net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2025__B _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2740__S _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2978__A2 _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[32\]_D u_arbiter.i_wb_cpu_rdt\[29\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1789__I0 _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2400_ _0415_ _0539_ _0562_ _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3380_ u_scanchain_local.data_out net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout102_I net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2331_ _0497_ _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2262_ _0423_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\] _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_78_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2193_ u_arbiter.i_wb_cpu_rdt\[16\] _0368_ _0323_ u_arbiter.i_wb_cpu_dbus_dat\[16\]
+ _0361_ u_arbiter.i_wb_cpu_dbus_dat\[17\] _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__2666__A1 u_cpu.cpu.immdec.imm19_12_20\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3128__CLK net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1949__B u_cpu.rf_ram.regzero vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2969__A2 _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2624__I u_cpu.cpu.csr_imm vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[23\]_D u_arbiter.i_wb_cpu_rdt\[20\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout15_I net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1977_ _1064_ net8 _1384_ _1234_ u_cpu.rf_ram.addr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_14_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2529_ _0677_ _0679_ _0680_ _0474_ _0477_ _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_121_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2409__A1 _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2409__B2 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[14\]_D u_arbiter.i_wb_cpu_rdt\[11\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2345__B1 _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2896__A1 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2709__I _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2880_ _0771_ _0946_ _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1900_ _1336_ _0020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1831_ _1036_ _1270_ _1272_ _1048_ _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_31_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1762_ _1032_ _1037_ _1205_ _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_1693_ _1122_ _1150_ _1151_ _1152_ u_arbiter.o_wb_cpu_adr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_143_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2887__A1 _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2314_ _0250_ u_arbiter.i_wb_cpu_rdt\[13\] _0481_ _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2245_ u_arbiter.i_wb_cpu_rdt\[11\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[11\]
+ _0248_ _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2639__A1 u_cpu.cpu.immdec.imm19_12_20\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2176_ u_arbiter.i_wb_cpu_dbus_dat\[12\] _0358_ _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1862__A2 _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2290__S _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2022__C _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2878__A1 _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1589__B _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2264__I _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1608__I _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2869__A1 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1771__C _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2030_ u_cpu.cpu.genblk1.align.ctrl_misal _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_43_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2097__A2 _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_63_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2932_ u_arbiter.i_wb_cpu_rdt\[28\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[12\]
+ _0979_ _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3210__D u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2863_ _0931_ _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2794_ u_cpu.cpu.ctrl.o_ibus_adr\[6\] _0885_ _0887_ u_cpu.cpu.ctrl.o_ibus_adr\[7\]
+ _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1814_ _1044_ _1243_ _1249_ u_cpu.cpu.genblk3.csr.mstatus_mie _1256_ _1257_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_1745_ u_arbiter.i_wb_cpu_dbus_adr\[29\] _1116_ _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2557__B1 _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1676_ u_arbiter.i_wb_cpu_dbus_adr\[14\] _1122_ _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1780__A1 _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2309__B1 _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout82_I net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2349__I _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2228_ _0401_ _0072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2159_ _0346_ _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2285__S _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1835__A2 u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2796__B1 _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1599__A1 _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2812__I _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1856__C _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2012__A2 _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2866__A4 _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2079__A2 _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1826__A2 u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2923__S _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_scanchain_local.scan_flop\[60\] u_scanchain_local.module_data_in\[59\] net146 u_arbiter.o_wb_cpu_adr\[22\]
+ net34 u_scanchain_local.module_data_in\[60\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__2003__A2 _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3200_ u_cpu.rf_ram_if.wdata0_r\[2\] net40 u_cpu.rf_ram_if.wdata0_r\[1\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[51\]_SE net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2169__I _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3131_ _0153_ net103 u_cpu.cpu.ctrl.o_ibus_adr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3205__D u_cpu.cpu.o_wdata0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3062_ _0087_ net55 u_cpu.cpu.decode.op22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2013_ _1231_ _0237_ _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2118__B _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2490__A2 _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2227__C1 _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2915_ _0972_ _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2846_ u_cpu.cpu.ctrl.o_ibus_adr\[28\] _0913_ _0915_ u_cpu.cpu.ctrl.o_ibus_adr\[29\]
+ _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_136_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2777_ net2 _0238_ _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1728_ u_arbiter.i_wb_cpu_dbus_adr\[25\] _1172_ _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1753__A1 u_arbiter.i_wb_cpu_dbus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1659_ _1124_ _1120_ _1125_ _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2233__A2 _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1992__A1 _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3011__CLK net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2472__A2 _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1777__B u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3161__CLK net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2700_ _0832_ _0113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2631_ _0500_ _0483_ _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_12_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2562_ _0476_ _0687_ _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2493_ u_cpu.cpu.immdec.imm24_20\[3\] _0640_ _0638_ _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3114_ _0139_ net118 u_arbiter.i_wb_cpu_dbus_adr\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3045_ _0070_ net93 u_arbiter.i_wb_cpu_dbus_dat\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout45_I net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2215__A2 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2362__I _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1974__A1 _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2829_ _0909_ _0165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1907__S net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2738__S _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3034__CLK net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3184__CLK net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2206__A2 _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout83 net84 net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout61 net62 net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_11_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout72 net85 net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout50 net59 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_122_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout94 net95 net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_31_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1965__A1 _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1616__I _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[23\] u_arbiter.i_wb_cpu_rdt\[20\] net128 u_arbiter.i_wb_cpu_dbus_dat\[17\]
+ net14 u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_81_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1993_ u_cpu.cpu.state.init_done _0219_ _0220_ _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_14_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2614_ _0730_ _0756_ _0758_ _0586_ _0101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2545_ _0420_ _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3057__CLK net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2476_ _0466_ _0500_ _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2558__S _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2133__A1 u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2684__A2 _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3028_ _0053_ net102 u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2436__A2 _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2675__A2 _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[33\]_CLK net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[48\]_CLK net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2330_ _0476_ _0496_ _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2261_ _0249_ _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2115__A1 _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2192_ _0376_ _0377_ _0060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2910__I0 u_arbiter.i_wb_cpu_rdt\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2666__A2 _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1874__B1 _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2905__I _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1976_ u_cpu.cpu.immdec.imm11_7\[1\] _1350_ net8 _1383_ _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_18_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2354__A1 _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2528_ u_arbiter.i_wb_cpu_rdt\[25\] u_arbiter.i_wb_cpu_rdt\[9\] _0590_ _0680_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1952__I1 _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2459_ _0482_ _0556_ _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2106__A1 u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2657__A2 _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2815__I _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2345__B2 _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2345__A1 _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2896__A2 _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[2\]_SE net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2820__A2 _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1830_ u_cpu.cpu.branch_op _1271_ _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__2584__A1 _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1761_ _1204_ u_cpu.cpu.bufreg.i_sh_signed _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1692_ u_arbiter.i_wb_cpu_dbus_adr\[17\] _1130_ _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2336__A1 _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2313_ _1078_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[13\] _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2887__A2 _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2244_ _0412_ _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2639__A2 _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2175_ _0363_ _0365_ _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2575__A1 _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1959_ _1372_ _0004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2575__B2 _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1915__S _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2878__A2 _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2545__I _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2566__A1 _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2869__A2 _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2931_ _0981_ _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1852__I0 _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2862_ _0513_ _0930_ _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2793_ _0888_ _0150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1813_ _1255_ _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2557__A1 _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1744_ u_cpu.cpu.ctrl.o_ibus_adr\[29\] _1191_ _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_50_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2557__B2 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1675_ _1111_ _1136_ _1137_ _1138_ u_arbiter.o_wb_cpu_adr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__2309__A1 _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2309__B2 _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1907__I1 u_cpu.rf_ram.data\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout75_I net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2227_ u_arbiter.i_wb_cpu_rdt\[27\] _0368_ _0390_ u_arbiter.i_wb_cpu_dbus_dat\[27\]
+ _0346_ u_arbiter.i_wb_cpu_dbus_dat\[28\] _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2158_ _0350_ _0353_ _0050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2089_ _1045_ _0287_ _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1599__A2 _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2548__A1 _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1619__I _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[53\] u_scanchain_local.module_data_in\[52\] net143 u_arbiter.o_wb_cpu_adr\[15\]
+ net29 u_scanchain_local.module_data_in\[53\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__2539__A1 _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1762__A2 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3130_ _0152_ net107 u_cpu.cpu.ctrl.o_ibus_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3061_ _0086_ net72 u_cpu.cpu.decode.op21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2012_ _1268_ _1273_ _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2227__B1 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2914_ u_arbiter.i_wb_cpu_rdt\[20\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[4\]
+ _0967_ _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2845_ _0918_ _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2776_ _0876_ _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1727_ u_cpu.cpu.ctrl.o_ibus_adr\[25\] _1178_ _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_144_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1753__A2 _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1658_ _1124_ _1120_ _1093_ _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2163__C1 _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1589_ _1066_ _1067_ _1023_ _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_6_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1992__A2 _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2941__A1 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2934__S _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2209__B1 _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout125_I net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2630_ _0516_ _0770_ _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_127_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2561_ _0537_ _0709_ _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_12_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2492_ u_cpu.cpu.immdec.imm24_20\[2\] _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3216__D u_cpu.rf_ram_if.wdata1_r\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3113_ _0138_ net117 u_arbiter.i_wb_cpu_dbus_adr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2160__A2 _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3044_ _0069_ net94 u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2129__B _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1671__A1 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2828_ _1160_ _0906_ _0908_ u_cpu.cpu.ctrl.o_ibus_adr\[21\] _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2759_ u_arbiter.i_wb_cpu_dbus_adr\[31\] _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1923__S _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout40 net42 net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA_u_scanchain_local.scan_flop\[41\]_SE net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout73 net78 net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout62 net86 net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_80_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout51 net54 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_11_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout95 net96 net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout84 net85 net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_35_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_scanchain_local.scan_flop\[16\] u_arbiter.i_wb_cpu_rdt\[13\] net130 u_arbiter.i_wb_cpu_dbus_dat\[10\]
+ net16 u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_93_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2693__A3 u_cpu.cpu.genblk3.csr.i_mtip vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1653__A1 u_arbiter.i_wb_cpu_dbus_adr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2850__B1 _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1992_ _1320_ _1266_ _0220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2613_ u_cpu.cpu.immdec.imm19_12_20\[1\] _0505_ _0757_ _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2544_ _0672_ _0692_ _0693_ _0676_ _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_130_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2475_ _0620_ _0630_ _0632_ _0533_ _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_141_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3027_ _0052_ net91 u_arbiter.i_wb_cpu_dbus_dat\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_97_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_109_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3001__CLK net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1580__B1 _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3151__CLK net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2832__B1 _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1635__A1 _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2060__A1 _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2260_ _0428_ _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2191_ u_arbiter.i_wb_cpu_rdt\[15\] _0364_ _0371_ u_arbiter.i_wb_cpu_dbus_dat\[15\]
+ _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1874__B2 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1874__A1 _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3024__CLK net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1975_ u_cpu.cpu.decode.op26 u_cpu.cpu.decode.co_ebreak _1341_ _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_14_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2051__A1 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2729__I1 u_arbiter.i_wb_cpu_dbus_adr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3174__CLK net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2527_ _0592_ _0503_ _0678_ _0529_ _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2458_ u_arbiter.i_wb_cpu_rdt\[26\] u_arbiter.i_wb_cpu_rdt\[10\] _0589_ _0616_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_130_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2106__A2 _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2368__I _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2389_ _0552_ _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_5_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1865__A1 _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1617__A1 u_arbiter.i_wb_cpu_dbus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2593__A2 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2345__A2 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[9\] u_arbiter.i_wb_cpu_rdt\[6\] net136 u_arbiter.i_wb_cpu_dbus_dat\[3\]
+ net21 u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_0_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1856__A1 _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1910__I _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3047__CLK net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2281__A1 _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1760_ u_arbiter.i_wb_cpu_dbus_we _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3197__CLK net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2584__A2 _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1691_ u_cpu.cpu.ctrl.o_ibus_adr\[17\] _1147_ _1145_ _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_7_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2336__A2 _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2312_ _0479_ _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2243_ _0411_ _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2174_ u_arbiter.i_wb_cpu_rdt\[10\] _0364_ _0348_ u_arbiter.i_wb_cpu_dbus_dat\[10\]
+ _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_66_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2916__I _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout20_I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1976__B net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2024__A1 _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1958_ u_cpu.rf_ram_if.rdata0\[5\] _1361_ _1057_ _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1889_ _0041_ _1322_ _1329_ _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2327__A2 _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2878__A3 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[32\]_CLK net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[47\]_CLK net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2263__A1 _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2015__A1 _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2566__A2 u_arbiter.i_wb_cpu_rdt\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2510__B _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_63_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2930_ u_arbiter.i_wb_cpu_rdt\[27\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[11\]
+ _0979_ _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_15_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2861_ _0218_ _0242_ _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2792_ _1100_ _0885_ _0887_ u_cpu.cpu.ctrl.o_ibus_adr\[6\] _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2404__C _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1812_ u_cpu.cpu.genblk3.csr.mcause3_0\[0\] _1250_ _1252_ _1254_ _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1743_ u_cpu.cpu.ctrl.o_ibus_adr\[28\] u_cpu.cpu.ctrl.o_ibus_adr\[27\] u_cpu.cpu.ctrl.o_ibus_adr\[26\]
+ _1182_ _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__2557__A2 _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3219__D u_cpu.cpu.o_wdata1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1674_ u_arbiter.i_wb_cpu_dbus_adr\[13\] _1130_ _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3212__CLK net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2226_ _0398_ _0394_ _0354_ _0399_ _0400_ _0071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout68_I net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2157_ u_arbiter.i_wb_cpu_dbus_dat\[5\] _0351_ _0352_ _0264_ _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1550__I _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2088_ _0293_ _0039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2796__A2 _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2548__A2 _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1926__S _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2757__S _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2484__A1 _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2236__A1 u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_scanchain_local.scan_flop\[46\] u_scanchain_local.module_data_in\[45\] net146 u_arbiter.o_wb_cpu_adr\[8\]
+ net34 u_scanchain_local.module_data_in\[46\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_10_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3060_ _0085_ net55 u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2011_ _1293_ _1280_ _0235_ _1287_ _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__2475__B2 _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2227__A1 u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2913_ _0971_ _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2844_ u_cpu.cpu.ctrl.o_ibus_adr\[27\] _0913_ _0915_ u_cpu.cpu.ctrl.o_ibus_adr\[28\]
+ _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_89_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2775_ _0875_ _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1726_ u_cpu.cpu.ctrl.o_ibus_adr\[24\] _1169_ _1170_ _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1657_ u_cpu.cpu.ctrl.o_ibus_adr\[10\] _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2950__A2 _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1545__I u_cpu.cpu.bufreg.lsb\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1588_ _1041_ _1044_ _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2163__C2 u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2163__B1 _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2209_ u_arbiter.i_wb_cpu_rdt\[21\] _0380_ _0351_ u_arbiter.i_wb_cpu_dbus_dat\[21\]
+ _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2466__A1 _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3189_ _0017_ net54 u_cpu.rf_ram.rdata\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2309__C _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2218__A1 u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3108__CLK net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[2\]_D net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2457__A1 u_cpu.cpu.decode.op26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2209__A1 u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout118_I net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2560_ _0620_ _0706_ _0708_ _0603_ _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_12_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2491_ _0601_ _0646_ _0090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3112_ _0137_ net120 u_arbiter.i_wb_cpu_dbus_adr\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3043_ _0068_ net97 u_arbiter.i_wb_cpu_dbus_dat\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2196__I _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2448__A1 _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2620__B2 _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2827_ _0878_ _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2758_ _0863_ _0140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1709_ u_arbiter.i_wb_cpu_dbus_adr\[21\] _1109_ _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2689_ u_cpu.cpu.immdec.imm31 _0489_ _0511_ _0823_ _0824_ _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_99_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2439__A1 _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout30 net36 net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout74 net78 net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout41 net42 net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3080__CLK net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout52 net54 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout63 net65 net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_70_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout96 net100 net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout85 net86 net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_11_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2678__A1 _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1653__A2 _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2850__B2 u_cpu.cpu.ctrl.o_ibus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1991_ _0218_ _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2612_ _0754_ _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2543_ _0545_ _0535_ _0491_ _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2474_ _0475_ _0631_ _0582_ _0621_ _0433_ _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__2669__A1 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout50_I net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3026_ _0051_ net101 u_arbiter.i_wb_cpu_dbus_dat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_u_scanchain_local.scan_flop\[26\]_D u_arbiter.i_wb_cpu_rdt\[23\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1883__A2 u_cpu.cpu.ctrl.i_iscomp vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[17\]_D u_arbiter.i_wb_cpu_rdt\[14\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2060__A2 _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2899__B2 _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2899__A1 _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2190_ u_arbiter.i_wb_cpu_dbus_dat\[16\] _0375_ _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1874__A2 _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1626__A2 _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1974_ _1069_ _1380_ _1381_ _1382_ u_cpu.rf_ram.addr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_14_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2423__B _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout98_I net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2526_ _0553_ _0533_ _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2457_ u_cpu.cpu.decode.op26 _0413_ _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1553__I _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2388_ _0424_ _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1865__A2 _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1617__A2 _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2384__I _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3009_ _0034_ net69 u_cpu.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2042__A2 u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2281__A2 _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1690_ _1147_ _1145_ u_cpu.cpu.ctrl.o_ibus_adr\[17\] _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_87_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1919__I0 u_cpu.rf_ram_if.wdata0_r\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout100_I net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[54\]_SE net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2311_ u_arbiter.i_wb_cpu_rdt\[14\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[14\]
+ _0416_ _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_48_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2242_ _0410_ _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2173_ _0338_ _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1847__A2 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xserv_0_160 io_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_90_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1976__C _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3141__CLK net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout13_I net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1548__I _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1957_ _1371_ _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1783__A1 _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1888_ _1327_ _1328_ _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2509_ _0414_ _0485_ _0491_ _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2263__A2 u_arbiter.i_wb_cpu_rdt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_123_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3014__CLK net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3164__CLK net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_fanout148_I net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2860_ _0246_ _0238_ _0928_ _0929_ _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_30_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1811_ _1231_ _1253_ _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2791_ _0879_ _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1742_ _1174_ _1189_ _1190_ u_arbiter.o_wb_cpu_adr\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1673_ u_cpu.cpu.ctrl.o_ibus_adr\[13\] _1133_ _1129_ _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_50_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2420__C _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2190__A1 u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2225_ u_arbiter.i_wb_cpu_rdt\[26\] _0318_ _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2927__I _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2156_ _0345_ _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2493__A2 _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2087_ _1072_ u_cpu.cpu.state.o_cnt_r\[2\] _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_59_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2989_ _0027_ net68 u_cpu.rf_ram_if.rreq_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3037__CLK net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2484__A2 _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2236__A2 _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1995__A1 _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2505__C _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_scanchain_local.scan_flop\[39\] u_scanchain_local.module_data_in\[38\] net137 u_arbiter.o_wb_cpu_adr\[1\]
+ net23 u_scanchain_local.module_data_in\[39\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_136_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2010_ _1293_ _1291_ _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2227__A2 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2912_ u_arbiter.i_wb_cpu_rdt\[19\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[3\]
+ _0967_ _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1986__A1 _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2843_ _0917_ _0171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2774_ _1231_ _0237_ net2 _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1725_ _1174_ _1176_ _1177_ u_arbiter.o_wb_cpu_adr\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1656_ u_arbiter.i_wb_cpu_dbus_adr\[10\] _1122_ _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_u_scanchain_local.scan_flop\[46\]_CLK net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2150__C _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1587_ _1047_ _1045_ _1050_ _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_59_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2163__A1 u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout80_I net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2208_ u_arbiter.i_wb_cpu_dbus_dat\[22\] _0352_ _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3188_ _0209_ net68 u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2139_ u_arbiter.i_wb_cpu_rdt\[3\] _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2218__A2 _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1977__B2 _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2154__A1 u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2457__A2 _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2209__A2 _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1968__A1 u_cpu.raddr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2490_ u_cpu.cpu.immdec.imm24_20\[2\] _0640_ _0645_ _0489_ _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2145__A1 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3111_ _0136_ net120 u_arbiter.i_wb_cpu_dbus_adr\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3042_ _0067_ net93 u_arbiter.i_wb_cpu_dbus_dat\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2426__B _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2826_ _0907_ _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2620__A2 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2757_ u_arbiter.i_wb_cpu_dbus_adr\[29\] u_arbiter.i_wb_cpu_dbus_adr\[30\] _0830_
+ _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1708_ u_cpu.cpu.ctrl.o_ibus_adr\[21\] _1163_ _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2688_ _0766_ _0719_ _0620_ _0530_ _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_133_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1639_ _1090_ _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_63_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2439__A2 _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout31 net32 net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout20 net38 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout42 net43 net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout53 net54 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout64 net65 net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout97 net98 net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout86 net125 net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout75 net77 net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_35_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2375__A1 _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2127__A1 _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2678__A2 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[5\]_SE net136 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2850__A2 _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1990_ u_cpu.cpu.state.o_cnt_r\[1\] _1281_ _1244_ u_cpu.cpu.state.o_cnt_r\[2\] _0218_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout130_I net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2611_ _0755_ _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2542_ _0487_ _0631_ _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2366__A1 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2473_ _0458_ _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2669__A2 _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3025_ _0050_ net101 u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_37_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout43_I net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2809_ _0897_ _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1580__A2 _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1950__S u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2832__A2 _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[21\] u_arbiter.i_wb_cpu_rdt\[18\] net127 u_arbiter.i_wb_cpu_dbus_dat\[15\]
+ net13 u_arbiter.i_wb_cpu_rdt\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_3_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1571__A2 _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2520__A1 _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2587__A1 _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1973_ u_cpu.cpu.immdec.imm11_7\[0\] _1341_ _1262_ _1380_ _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_53_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2525_ _0533_ _0674_ _0676_ _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1562__A2 u_cpu.cpu.decode.op26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2456_ _1245_ _0587_ _0614_ _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_64_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3070__CLK net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2387_ _0475_ _0543_ _0544_ _0467_ _0550_ _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3008_ _0033_ net79 u_cpu.cpu.state.o_cnt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2578__A1 _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2524__B _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xu_scanchain_local.scan_flop\[69\] u_scanchain_local.module_data_in\[68\] net147 u_arbiter.o_wb_cpu_adr\[31\]
+ net31 u_scanchain_local.module_data_in\[69\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__2569__A1 _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3093__CLK net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1919__I1 u_cpu.rf_ram_if.wdata1_r\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2310_ _0224_ _0413_ _0451_ _0478_ _0077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_3_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2241_ net12 _1073_ _0409_ _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2172_ u_arbiter.i_wb_cpu_dbus_dat\[11\] _0358_ _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1956_ u_cpu.rf_ram_if.rdata0\[4\] _1359_ u_cpu.rf_ram_if.rtrig0 _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2980__A1 _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1887_ _1265_ _1321_ _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2193__C1 _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2508_ _0642_ _0659_ _0660_ _0661_ _0092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_130_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2439_ _0487_ _0544_ _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2609__B _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2239__B1 _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1810_ _1040_ u_cpu.cpu.decode.co_ebreak _1043_ _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_15_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[21\]_SE net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2790_ _0886_ _0149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1741_ u_arbiter.i_wb_cpu_dbus_adr\[28\] _1116_ _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1672_ _1133_ _1129_ u_cpu.cpu.ctrl.o_ibus_adr\[13\] _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_139_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2190__A2 _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2224_ u_arbiter.i_wb_cpu_dbus_dat\[27\] _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_61_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2155_ _0322_ _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2086_ _0247_ _1323_ _0038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_4_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2988_ _0269_ _1019_ _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1939_ _1360_ _0009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2953__A1 _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1692__A1 u_arbiter.i_wb_cpu_dbus_adr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[44\]_SE net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1995__A2 _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2172__A2 _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3131__CLK net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2911_ _0970_ _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_cpu.rf_ram.RAM0_A[7] u_cpu.rf_ram.addr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1986__A2 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2842_ _1181_ _0913_ _0915_ u_cpu.cpu.ctrl.o_ibus_adr\[27\] _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_32_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2773_ _0216_ _0870_ _0874_ _0144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1724_ u_arbiter.i_wb_cpu_dbus_adr\[24\] _1172_ _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2999__CLK net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1655_ _1090_ _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1586_ u_cpu.cpu.immdec.imm19_12_20\[6\] _1027_ _1055_ u_cpu.cpu.immdec.imm24_20\[2\]
+ _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__2163__A2 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout73_I net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2207_ _0386_ _0387_ _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2466__A3 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3187_ _0208_ net74 u_cpu.cpu.ctrl.i_iscomp vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[67\]_SE net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2138_ _0336_ _0047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2069_ _1244_ u_cpu.cpu.state.o_cnt\[2\] _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_50_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1977__A2 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2622__B _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3004__CLK net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2154__A2 _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2090__A1 _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[51\] u_scanchain_local.module_data_in\[50\] net141 u_arbiter.o_wb_cpu_adr\[13\]
+ net28 u_scanchain_local.module_data_in\[51\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_51_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.out_flop u_scanchain_local.module_data_in\[69\] net31 u_scanchain_local.data_out_i
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XANTENNA__2145__A2 _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3110_ _0135_ net120 u_arbiter.i_wb_cpu_dbus_adr\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3041_ _0066_ net97 u_arbiter.i_wb_cpu_dbus_dat\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3027__CLK net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2825_ u_cpu.cpu.ctrl.o_ibus_adr\[19\] _0906_ _0901_ _1160_ _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_32_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2442__B _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2756_ _0862_ _0139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1707_ _1160_ _1157_ _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2687_ u_arbiter.i_wb_cpu_rdt\[31\] u_arbiter.i_wb_cpu_rdt\[15\] _1083_ _0823_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1638_ u_cpu.cpu.ctrl.o_ibus_adr\[7\] _1105_ _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_132_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1569_ u_cpu.cpu.decode.opcode\[2\] _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_24_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout21 net22 net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout10 net11 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_70_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout32 net35 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_35_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout43 net44 net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__2072__A1 _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout65 net66 net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout54 net58 net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout98 net99 net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout87 net90 net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_12
Xfanout76 net77 net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_109_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2375__A2 _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[45\]_CLK net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2063__A1 _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout123_I net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2610_ _0754_ _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2541_ _0637_ _0691_ _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2472_ _0622_ _0485_ _0544_ _0546_ _0629_ _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_130_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1629__A1 u_cpu.cpu.genblk1.align.ctrl_misal vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3024_ _0049_ net101 u_arbiter.i_wb_cpu_dbus_dat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1644__A4 _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout36_I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1567__I _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2808_ _1133_ _0892_ _0894_ u_cpu.cpu.ctrl.o_ibus_adr\[13\] _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2739_ _0853_ _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2357__A2 u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2109__A2 u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2398__I _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2668__I0 u_arbiter.i_wb_cpu_rdt\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2045__A1 _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2596__A2 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_scanchain_local.scan_flop\[14\] u_arbiter.i_wb_cpu_rdt\[11\] net134 u_arbiter.i_wb_cpu_dbus_dat\[8\]
+ net20 u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_46_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2808__B1 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2284__A1 _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1972_ _1041_ _1234_ _1350_ _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_18_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2339__A2 _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2524_ _0553_ _0675_ _0624_ _0575_ _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_2455_ _0588_ _0602_ _0613_ _0498_ _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3215__CLK net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2386_ _0525_ _0547_ _0549_ _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_57_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3007_ _0032_ net80 u_cpu.cpu.state.stage_two_req vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2027__A1 _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2578__A2 _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2266__A1 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2524__C _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2569__A2 _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2240_ _0251_ u_arbiter.i_wb_cpu_ibus_adr\[1\] _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2171_ _0362_ _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_47_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_cpu.rf_ram.RAM0_D[7] u_cpu.rf_ram.i_wdata\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1955_ _1370_ _0002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1886_ _1325_ _1326_ _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_128_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2193__B1 _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2193__C2 u_arbiter.i_wb_cpu_dbus_dat\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2507_ u_cpu.cpu.immdec.imm24_20\[3\] _0642_ _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2438_ _0507_ _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2496__A1 _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2369_ _0502_ _0457_ _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1956__S u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2420__B2 _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2420__A1 _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2184__B1 _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[7\] u_arbiter.i_wb_cpu_rdt\[4\] net137 u_arbiter.i_wb_cpu_dbus_dat\[1\]
+ net21 u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_43_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2239__B2 _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2535__B _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1740_ u_cpu.cpu.ctrl.o_ibus_adr\[28\] _1188_ _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2411__A1 _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1671_ _1132_ _1134_ _1135_ u_arbiter.o_wb_cpu_adr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2223_ u_arbiter.i_wb_cpu_dbus_dat\[26\] _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2478__A1 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2154_ u_arbiter.i_wb_cpu_rdt\[5\] _0339_ _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2085_ _0292_ _0037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2650__A1 _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1989__B1 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2987_ _0255_ _1018_ _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2402__A1 _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1938_ u_cpu.rf_ram_if.rdata1\[3\] _1359_ _1355_ _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1869_ _1310_ _1272_ _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2469__A1 _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1692__A2 _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2157__B1 _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[5\]_D u_arbiter.i_wb_cpu_rdt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2910_ u_arbiter.i_wb_cpu_rdt\[18\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[2\]
+ _0967_ _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_44_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2632__A1 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_cpu.rf_ram.RAM0_A[6] u_cpu.rf_ram.addr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2841_ _0916_ _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_32_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2772_ _0870_ _0873_ _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_89_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1723_ u_cpu.cpu.ctrl.o_ibus_adr\[24\] _1175_ _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_89_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1654_ _1111_ _1118_ _1120_ _1121_ u_arbiter.o_wb_cpu_adr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1585_ u_cpu.cpu.immdec.imm19_12_20\[5\] _1057_ _1063_ _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_99_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2206_ u_arbiter.i_wb_cpu_rdt\[20\] _0380_ _0351_ u_arbiter.i_wb_cpu_dbus_dat\[20\]
+ _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_26_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout66_I net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3186_ _0207_ net71 u_cpu.cpu.genblk3.csr.mstatus_mie vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2320__B1 _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1674__A2 _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2137_ u_arbiter.i_wb_cpu_rdt\[2\] _0318_ _0335_ _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2871__B2 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2068_ _1244_ u_cpu.cpu.state.o_cnt\[2\] _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2623__B2 _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2387__B1 _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1665__A2 _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2862__A1 _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2614__A1 _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2614__B2 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[44\] u_scanchain_local.module_data_in\[43\] net147 u_arbiter.o_wb_cpu_adr\[6\]
+ net31 u_scanchain_local.module_data_in\[44\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_138_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3040_ _0065_ net99 u_arbiter.i_wb_cpu_dbus_dat\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1656__A2 _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2853__A1 _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[38\]_D u_scanchain_local.module_data_in\[37\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2081__A2 _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2824_ _0875_ _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2755_ u_arbiter.i_wb_cpu_dbus_adr\[28\] u_arbiter.i_wb_cpu_dbus_adr\[29\] _0830_
+ _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1706_ _1132_ _1161_ _1162_ u_arbiter.o_wb_cpu_adr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2686_ _0781_ _0818_ _0821_ _0822_ _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1637_ _1104_ _1106_ _1107_ u_arbiter.o_wb_cpu_adr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[34\]_SE net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1568_ u_cpu.cpu.genblk3.csr.o_new_irq _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_28_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3169_ _0190_ net88 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[29\]_D u_arbiter.i_wb_cpu_rdt\[26\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout22 net26 net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout11 _0026_ net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout33 net34 net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2633__B _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2072__A2 _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout44 net126 net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout55 net56 net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout99 net100 net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
Xfanout88 net90 net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout77 net78 net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_35_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout66 net72 net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_127_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3121__CLK net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1583__A1 u_cpu.cpu.decode.op26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2780__B1 _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2989__CLK net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2527__C _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2543__B _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1810__A2 u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout116_I net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2540_ u_cpu.cpu.immdec.imm30_25\[1\] _0688_ _0690_ u_cpu.cpu.immdec.imm30_25\[2\]
+ _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_142_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2471_ _0626_ _0628_ _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__1574__A1 _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1877__A2 _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3023_ _0048_ net104 u_arbiter.i_wb_cpu_dbus_dat\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1629__A2 u_cpu.cpu.ctrl.o_ibus_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3144__CLK net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout29_I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2054__A2 _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2807_ _0896_ _0156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_34_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2738_ u_arbiter.i_wb_cpu_dbus_adr\[20\] u_arbiter.i_wb_cpu_dbus_adr\[21\] _0849_
+ _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1565__A1 _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2669_ _0631_ _0484_ _0576_ _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2514__B1 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2668__I1 u_arbiter.i_wb_cpu_rdt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2293__A2 u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1758__I _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3017__CLK net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2284__A2 u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1971_ _1202_ _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_18_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2523_ _0593_ _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2454_ _0603_ _0610_ _0611_ _0612_ _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_116_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2385_ _0548_ _0482_ _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput1 io_in[0] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__2275__A2 _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3006_ _0006_ net45 u_cpu.rf_ram_if.rdata0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[44\]_CLK net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1710__A1 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[59\]_CLK net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2018__A2 _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2112__I _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2170_ u_arbiter.i_wb_cpu_rdt\[9\] _0321_ _0323_ u_arbiter.i_wb_cpu_dbus_dat\[9\]
+ _0361_ u_arbiter.i_wb_cpu_dbus_dat\[10\] _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_4_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_cpu.rf_ram.RAM0_D[6] u_cpu.rf_ram.i_wdata\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1954_ u_cpu.rf_ram_if.rdata0\[3\] _1357_ u_cpu.rf_ram_if.rtrig0 _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1885_ _1071_ u_cpu.cpu.ctrl.pc_plus_4_cy_r _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_128_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2193__A1 u_arbiter.i_wb_cpu_rdt\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2193__B2 u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout96_I net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2506_ u_cpu.cpu.immdec.imm24_20\[4\] _0568_ _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2437_ _0592_ _0595_ _0596_ _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2368_ _0429_ _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2299_ _0466_ _0467_ _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2420__A2 _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2184__A1 u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2487__A2 _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2239__A2 _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1670_ u_arbiter.i_wb_cpu_dbus_adr\[12\] _1109_ _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2222_ _0397_ _0070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2153_ _0347_ _0349_ _0049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2084_ _0282_ _1281_ _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1989__A1 _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2650__A2 _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout11_I _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2986_ _1016_ _1017_ _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2402__A2 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1937_ _1353_ _0020_ _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1868_ _1030_ _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1799_ _1236_ _1241_ _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_40_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2157__B2 _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2157__A1 u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_u_scanchain_local.scan_flop\[8\]_SE net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1683__A3 _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_cpu.rf_ram.RAM0_A[5] u_cpu.rf_ram.addr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2840_ u_cpu.cpu.ctrl.o_ibus_adr\[25\] _0913_ _0915_ _1181_ _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2632__A2 _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_106_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2771_ _0868_ _0872_ _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2396__A1 _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1722_ _1169_ _1170_ _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1653_ u_arbiter.i_wb_cpu_dbus_adr\[9\] _1116_ _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1584_ _1024_ _1038_ _1061_ _1062_ _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_85_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2205_ u_arbiter.i_wb_cpu_dbus_dat\[21\] _0375_ _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2320__A1 _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2320__B2 _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3185_ _0206_ net68 u_cpu.cpu.genblk3.csr.mie_mtie vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2136_ _0331_ _0333_ _0267_ _0334_ _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA_fanout59_I net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2456__B _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2067_ _0279_ _0032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2623__A2 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2969_ u_cpu.cpu.genblk3.csr.mstatus_mpie _1038_ _1234_ _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2387__A1 _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2387__B2 _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2934__I0 u_arbiter.i_wb_cpu_rdt\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3050__CLK net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2862__A2 _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2614__A2 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[37\] u_scanchain_local.module_data_in\[36\] net137 u_arbiter.i_wb_cpu_dbus_dat\[31\]
+ net24 u_scanchain_local.module_data_in\[37\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_49_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2925__I0 u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2550__A1 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2302__A1 _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2853__A2 _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2605__A2 _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2823_ _0905_ _0163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_56_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2754_ _0861_ _0138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2369__A1 _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1705_ u_arbiter.i_wb_cpu_dbus_adr\[20\] _1109_ _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2685_ u_cpu.cpu.immdec.imm19_12_20\[8\] _0755_ _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1636_ u_arbiter.i_wb_cpu_dbus_adr\[6\] _1091_ _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3073__CLK net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1567_ _1045_ _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2030__I u_cpu.cpu.genblk1.align.ctrl_misal vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3168_ _0189_ net88 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2119_ net12 _1089_ _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_55_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3099_ _0124_ net97 u_arbiter.i_wb_cpu_dbus_adr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout12 u_arbiter.i_wb_cpu_ack net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout34 net35 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout23 net24 net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout45 net46 net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout56 net57 net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout89 net90 net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout78 net84 net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout67 net71 net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_11_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1958__I1 _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2780__A1 _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2780__B2 u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1583__A2 u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2532__A1 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3096__CLK net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout109_I net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2470_ _0438_ _0464_ _0627_ _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1574__A2 _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3022_ _0047_ net105 u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2453__C _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2806_ u_cpu.cpu.ctrl.o_ibus_adr\[11\] _0892_ _0894_ _1133_ _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2737_ _0852_ _0130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2668_ u_arbiter.i_wb_cpu_rdt\[18\] u_arbiter.i_wb_cpu_rdt\[2\] _0590_ _0806_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1565__A2 _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2762__A1 u_cpu.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1619_ _1089_ _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2599_ _0740_ _0741_ _0742_ _0744_ _0554_ _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2514__A1 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1774__I u_cpu.cpu.immdec.imm11_7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2505__A1 _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2808__A2 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1970_ _1379_ u_cpu.rf_ram.addr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_18_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[24\]_SE net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2441__B1 _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1547__A2 _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2522_ _0475_ _0673_ _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2453_ _0579_ _0545_ _0548_ _0602_ _0583_ _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2384_ _0506_ _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput2 io_in[1] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3111__CLK net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3005_ _0005_ net45 u_cpu.rf_ram_if.rdata0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1594__I u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2639__B _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[47\]_SE net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2974__A1 _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3134__CLK net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2549__B _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1701__A2 _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_cpu.rf_ram.RAM0_D[5] u_cpu.rf_ram.i_wdata\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2662__B1 _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xserv_0_153 io_oeb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_94_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1953_ _1369_ _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1884_ _1323_ u_cpu.cpu.ctrl.i_iscomp _1250_ _1324_ _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__2965__A1 _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2193__A2 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2505_ _0474_ _0649_ _0658_ _0477_ _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2436_ _0491_ _0486_ _0580_ _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_102_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1940__A2 _0021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout89_I net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2367_ _1209_ _0515_ _0532_ _0080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2740__I1 u_arbiter.i_wb_cpu_dbus_adr\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2298_ _0459_ _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3007__CLK net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3157__CLK net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2184__A2 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2495__I0 u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_106_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[67\] u_scanchain_local.module_data_in\[66\] net147 u_arbiter.o_wb_cpu_adr\[29\]
+ net31 u_scanchain_local.module_data_in\[67\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_15_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2221_ u_arbiter.i_wb_cpu_rdt\[25\] _0368_ _0390_ u_arbiter.i_wb_cpu_dbus_dat\[25\]
+ _0361_ u_arbiter.i_wb_cpu_dbus_dat\[26\] _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_87_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2152_ u_arbiter.i_wb_cpu_rdt\[4\] _0339_ _0348_ u_arbiter.i_wb_cpu_dbus_dat\[4\]
+ _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2083_ _0288_ _0291_ _0036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1989__A2 _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[43\]_CLK net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2985_ _0271_ u_cpu.rf_ram_if.rcnt\[1\] _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1936_ _1358_ _0008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1610__A1 _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1867_ _1289_ _1308_ _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_u_scanchain_local.scan_flop\[58\]_CLK net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1798_ _1237_ _1239_ _1240_ _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2166__A2 _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2419_ _0578_ _0579_ _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2636__C _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1601__A1 u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2157__A2 _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_cpu.rf_ram.RAM0_A[4] u_cpu.rf_ram.addr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1840__A1 _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2770_ u_arbiter.i_wb_cpu_dbus_adr\[2\] _0243_ _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout139_I net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1721_ _1093_ _1174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1652_ _1119_ _1112_ _1113_ _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_144_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2788__I _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2148__A2 _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1583_ u_cpu.cpu.decode.op26 u_cpu.cpu.decode.co_ebreak _1034_ _1042_ _1062_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_140_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2204_ _0384_ _0385_ _0064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3184_ _0205_ net67 u_cpu.cpu.genblk3.csr.mstatus_mpie vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2135_ u_arbiter.i_wb_cpu_dbus_dat\[2\] _0327_ _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2320__A2 _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2066_ _0246_ _0278_ _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2028__I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2084__A1 _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2968_ _0922_ _1249_ _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2387__A2 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1919_ u_cpu.rf_ram_if.wdata0_r\[4\] u_cpu.rf_ram_if.wdata1_r\[4\] _1342_ _1347_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2899_ _1389_ _0932_ _0963_ _0669_ _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2698__I _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2075__A1 _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1586__B1 _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2302__A2 _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2066__A1 _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2822_ u_cpu.cpu.ctrl.o_ibus_adr\[18\] _0899_ _0901_ u_cpu.cpu.ctrl.o_ibus_adr\[19\]
+ _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2753_ u_arbiter.i_wb_cpu_dbus_adr\[27\] u_arbiter.i_wb_cpu_dbus_adr\[28\] _0830_
+ _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2369__A2 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1704_ _1160_ _1157_ _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2512__S _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1577__B1 _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2684_ _1266_ _0732_ _0820_ _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1635_ _1075_ _1105_ _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1566_ u_cpu.cpu.state.genblk1.misalign_trap_sync_r _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_28_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout71_I net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3167_ _0188_ net88 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3098_ _0123_ net97 u_arbiter.i_wb_cpu_dbus_adr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2118_ net39 _0317_ _0318_ _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2049_ net12 _1088_ _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout13 net14 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout35 net36 net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout24 net25 net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1597__I _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1804__A1 _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout46 net50 net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout79 net80 net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout68 net70 net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout57 net58 net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_109_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1970__I _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3021_ _0046_ net101 u_arbiter.i_wb_cpu_dbus_dat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2039__A1 _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2306__I _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2805_ _0895_ _0155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3040__CLK net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2736_ u_arbiter.i_wb_cpu_dbus_adr\[19\] u_arbiter.i_wb_cpu_dbus_adr\[20\] _0849_
+ _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2762__A2 _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2667_ _0781_ _0803_ _0804_ _0805_ _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1618_ _1085_ _1087_ _1092_ u_arbiter.o_wb_cpu_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2598_ _0621_ _0519_ _0743_ _0579_ _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3190__CLK net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2514__A2 _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1880__I _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1549_ u_cpu.cpu.csr_d_sel _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_68_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3219_ u_cpu.cpu.o_wdata1 net56 u_cpu.rf_ram_if.wdata1_r\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1876__I1 u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2450__A1 _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2450__B2 _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2505__A2 _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2269__A1 _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3063__CLK net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2441__A1 _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout121_I net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2521_ _0495_ _0672_ _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2452_ _0441_ _0582_ _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2383_ _0545_ _0546_ _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3004_ _0004_ net51 u_cpu.rf_ram_if.rdata0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput3 io_in[2] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_92_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2680__A1 _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout34_I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2036__I _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2719_ _0842_ _0122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2499__A1 _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3086__CLK net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2671__A1 _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2423__A1 _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2974__A2 _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2187__B1 _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[12\] u_arbiter.i_wb_cpu_rdt\[9\] net135 u_arbiter.i_wb_cpu_dbus_dat\[6\]
+ net21 u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_4_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_cpu.rf_ram.RAM0_D[4] u_cpu.rf_ram.i_wdata\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2662__A1 _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xserv_0_154 io_oeb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2662__B2 _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2414__A1 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1952_ u_cpu.rf_ram_if.rdata0\[2\] _1354_ u_cpu.rf_ram_if.rtrig0 _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_15_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1883_ u_cpu.cpu.state.o_cnt_r\[2\] u_cpu.cpu.ctrl.i_iscomp _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2504_ _0583_ _0653_ _0655_ _0657_ _0496_ _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_2435_ _0486_ _0594_ _0575_ _0470_ _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_29_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2366_ _0517_ _0527_ _0531_ _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2297_ _0446_ _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2405__A1 _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2956__A2 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[10\]_D u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2892__A1 _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2644__A1 _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2495__I1 u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3101__CLK net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[8\]_D u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2220_ _0395_ _0396_ _0069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2151_ _0322_ _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_94_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2082_ _0282_ _0219_ _0290_ _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_59_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2984_ _1020_ _1022_ _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1935_ u_cpu.rf_ram_if.rdata1\[2\] _1357_ _1355_ _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1866_ _1258_ _1029_ u_cpu.cpu.alu.cmp_r _1307_ _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_1797_ _1237_ u_cpu.cpu.csr_imm _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[37\]_SE net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2418_ _0493_ _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2874__A1 _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2349_ _0514_ _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2626__A1 _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1601__A2 _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xu_scanchain_local.scan_flop\[5\] u_arbiter.i_wb_cpu_rdt\[2\] net136 u_arbiter.i_wb_cpu_dbus_sel\[3\]
+ net22 u_arbiter.i_wb_cpu_rdt\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2865__A1 _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2865__B2 _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2617__B2 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_cpu.rf_ram.RAM0_A[3] u_cpu.rf_ram.addr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1840__A2 _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_89_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1720_ _1132_ _1171_ _1173_ u_arbiter.o_wb_cpu_adr\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1651_ u_cpu.cpu.ctrl.o_ibus_adr\[9\] _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1582_ u_cpu.cpu.immdec.imm24_20\[1\] _1053_ _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2203_ u_arbiter.i_wb_cpu_rdt\[19\] _0380_ _0351_ u_arbiter.i_wb_cpu_dbus_dat\[19\]
+ _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3183_ _0204_ net67 u_cpu.cpu.genblk3.csr.mcause31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2134_ _0313_ _0332_ _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2065_ _0277_ _0257_ _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3147__CLK net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2084__A2 _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2967_ _0922_ _1260_ _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_120_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1918_ _1346_ u_cpu.rf_ram.i_wdata\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2898_ _0961_ _0962_ _0931_ _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2792__B1 _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1849_ u_cpu.cpu.mem_bytecnt\[1\] _1290_ _1224_ _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_2_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1586__A1 u_cpu.cpu.immdec.imm19_12_20\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[42\]_CLK net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2821_ _0904_ _0162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2752_ _0860_ _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1703_ u_cpu.cpu.ctrl.o_ibus_adr\[20\] _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2683_ _0530_ _0819_ _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1634_ u_cpu.cpu.ctrl.o_ibus_adr\[6\] _1100_ _1101_ _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_132_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1565_ _1039_ _1041_ _1043_ _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_28_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3166_ _0187_ net87 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout64_I net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3097_ _0122_ net97 u_arbiter.i_wb_cpu_dbus_adr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2117_ _0266_ _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2057__A2 _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2483__B _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2048_ _1258_ _1029_ _0264_ _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout14 net15 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout36 net37 net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout25 net26 net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout47 net49 net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_11_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout69 net70 net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout58 net59 net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__2703__S _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1788__I _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2048__A2 _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1559__A1 _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[42\] u_scanchain_local.module_data_in\[41\] net138 u_arbiter.o_wb_cpu_adr\[4\]
+ net23 u_scanchain_local.module_data_in\[42\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_6_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2568__B _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3020_ _0045_ net101 u_arbiter.i_wb_cpu_dbus_dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1899__S _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2804_ _1124_ _0892_ _0894_ u_cpu.cpu.ctrl.o_ibus_adr\[11\] _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2735_ _0851_ _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2666_ u_cpu.cpu.immdec.imm19_12_20\[6\] _0755_ _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1617_ u_arbiter.i_wb_cpu_dbus_adr\[2\] _1091_ _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2597_ _0740_ _0502_ _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2478__B _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1548_ _1023_ _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_80_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3218_ u_cpu.rf_ram_if.wdata1_r\[7\] net47 u_cpu.rf_ram_if.wdata1_r\[6\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3149_ _0171_ net117 u_cpu.cpu.ctrl.o_ibus_adr\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1876__I2 u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2202__A2 _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1713__A1 u_arbiter.i_wb_cpu_dbus_adr\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2269__A2 u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3208__CLK net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2441__A2 _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout114_I net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2520_ _0467_ _0464_ _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2451_ _0609_ _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1981__I _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2382_ u_arbiter.i_wb_cpu_rdt\[5\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\] _1080_
+ _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3003_ _0003_ net53 u_cpu.rf_ram_if.rdata0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput4 io_in[3] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_80_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2680__A2 _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2317__I _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout27_I net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2718_ u_arbiter.i_wb_cpu_dbus_adr\[11\] u_arbiter.i_wb_cpu_dbus_adr\[12\] _0837_
+ _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2649_ _0444_ _0773_ _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2743__I0 u_arbiter.i_wb_cpu_dbus_adr\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2671__A2 _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2423__A2 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2187__A1 u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_cpu.rf_ram.RAM0_D[3] u_cpu.rf_ram.i_wdata\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3030__CLK net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2111__A1 _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2662__A2 _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xserv_0_155 io_oeb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__3180__CLK net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2414__A2 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1951_ _1368_ _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1882_ u_cpu.cpu.state.o_cnt_r\[1\] _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_30_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2503_ _0546_ _0557_ _0656_ _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2434_ _0502_ _0593_ _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2725__I0 u_arbiter.i_wb_cpu_dbus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2365_ _0491_ _0528_ _0438_ _0529_ _0530_ _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_9_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2350__A1 _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2296_ _0460_ _0464_ _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__2102__A1 _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_75_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3053__CLK net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2877__C1 _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2644__A2 _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2332__A1 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2150_ u_arbiter.i_wb_cpu_dbus_dat\[5\] _0317_ _0260_ _0344_ _0346_ _0347_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2081_ _0289_ _0269_ _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2983_ _1015_ _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1934_ _1353_ _0019_ _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1865_ _1281_ _1247_ _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1796_ _1238_ _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3076__CLK net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout94_I net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2571__A1 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2417_ _0480_ _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2323__A1 _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2874__A2 _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2348_ _0513_ _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2279_ _0446_ _0447_ _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1921__I1 u_cpu.rf_ram_if.wdata1_r\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2626__A2 _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2562__A1 _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2617__A2 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_u_cpu.rf_ram.RAM0_A[2] u_cpu.rf_ram.addr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3099__CLK net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1650_ u_cpu.cpu.ctrl.o_ibus_adr\[9\] _1115_ _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2928__I0 u_arbiter.i_wb_cpu_rdt\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1581_ _1056_ _1058_ _1059_ _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_26_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2202_ u_arbiter.i_wb_cpu_dbus_dat\[20\] _0375_ _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3182_ _0203_ net67 u_cpu.cpu.genblk3.csr.mcause3_0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2133_ u_arbiter.i_wb_cpu_dbus_dat\[2\] _1317_ net39 _0314_ _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1903__I1 u_cpu.rf_ram.data\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2064_ _1217_ _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2966_ _1002_ _1004_ _1005_ _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_33_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1917_ u_cpu.rf_ram_if.wdata0_r\[3\] u_cpu.rf_ram_if.wdata1_r\[3\] _1342_ _1346_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2897_ _0412_ _0562_ _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1848_ u_cpu.cpu.state.o_cnt\[2\] u_cpu.cpu.mem_bytecnt\[0\] _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2919__I0 u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1779_ u_cpu.cpu.bufreg2.i_cnt_done u_cpu.cpu.immdec.imm31 _1222_ _1223_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[11\]_SI u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1586__A2 _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2535__A1 _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[27\]_SE net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2820_ u_cpu.cpu.ctrl.o_ibus_adr\[17\] _0899_ _0901_ u_cpu.cpu.ctrl.o_ibus_adr\[18\]
+ _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_fanout144_I net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2751_ u_arbiter.i_wb_cpu_dbus_adr\[26\] u_arbiter.i_wb_cpu_dbus_adr\[27\] _0855_
+ _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1702_ _1122_ _1157_ _1158_ _1159_ u_arbiter.o_wb_cpu_adr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__2774__A1 _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1577__A2 _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2682_ _1033_ u_cpu.cpu.immdec.imm24_20\[0\] _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1633_ _1100_ _1101_ u_cpu.cpu.ctrl.o_ibus_adr\[6\] _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2526__A1 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1564_ _1034_ _1042_ _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3114__CLK net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3165_ _0186_ net87 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3096_ _0121_ net111 u_arbiter.i_wb_cpu_dbus_adr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2116_ _0258_ _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_fanout57_I net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2047_ _0258_ _0261_ _0263_ _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_39_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout15 net19 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout26 net37 net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout37 net38 net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__1804__A3 u_cpu.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout48 net49 net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout59 net62 net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_2949_ u_cpu.cpu.genblk3.csr.mcause3_0\[3\] _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2765__B2 _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2004__B _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1843__B u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2048__A3 _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2453__B1 _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2508__A1 _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_scanchain_local.scan_flop\[35\] u_scanchain_local.module_data_in\[34\] net144 u_arbiter.i_wb_cpu_dbus_dat\[29\]
+ net30 u_scanchain_local.module_data_in\[35\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2568__C _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2584__B _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2803_ _0879_ _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2734_ u_arbiter.i_wb_cpu_dbus_adr\[18\] u_arbiter.i_wb_cpu_dbus_adr\[19\] _0849_
+ _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2665_ u_cpu.cpu.immdec.imm19_12_20\[7\] _0568_ _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1616_ _1090_ _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2596_ _0425_ _0582_ _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1547_ _1025_ _1026_ u_arbiter.i_wb_cpu_dbus_sel\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3217_ u_cpu.rf_ram_if.wdata1_r\[6\] net44 u_cpu.rf_ram_if.wdata1_r\[5\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3148_ _0170_ net117 u_cpu.cpu.ctrl.o_ibus_adr\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1876__I3 u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3079_ _0104_ net57 u_cpu.cpu.immdec.imm19_12_20\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2714__S _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[41\]_CLK net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[56\]_CLK net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2669__B _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1713__A2 _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout107_I net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2450_ _0605_ _0606_ _0607_ _0608_ _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_114_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2901__A1 _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1704__A2 _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2381_ u_arbiter.i_wb_cpu_rdt\[6\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[6\] _1080_
+ _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xinput5 io_in[4] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3002_ _0002_ net63 u_cpu.rf_ram_if.rdata0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2968__A1 _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1658__B _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2333__I _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2717_ _0841_ _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2648_ _0462_ _0741_ _0785_ _0787_ _0554_ _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2579_ _0695_ _0485_ _0718_ _0725_ _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2259__I0 u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2671__C _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2187__A2 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2431__I0 u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_cpu.rf_ram.RAM0_D[2] u_cpu.rf_ram.i_wdata\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2418__I _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xserv_0_156 io_oeb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1950_ u_cpu.rf_ram_if.rdata0\[1\] _1367_ u_cpu.rf_ram_if.rtrig0 _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1881_ _1237_ _1319_ _1320_ _1321_ _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_70_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2502_ _0471_ _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2433_ _0500_ _0482_ _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2364_ _0411_ _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2350__A2 _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2295_ _0463_ _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2810__B1 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1613__A1 _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1835__C u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2992__CLK net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2341__A2 _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2877__C2 _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2877__B1 _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[60\]_SE net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2801__B1 _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2332__A2 _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2080_ u_cpu.rf_ram_if.rgnt _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_4_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1987__I _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2982_ _0282_ u_cpu.rf_ram_if.rreq_r _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1933_ _1356_ _0007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1864_ _1237_ _1303_ _1304_ _1305_ _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__2611__I _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1795_ _1207_ _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2416_ _0533_ _0574_ _0576_ _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_fanout87_I net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2323__A2 _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2259__S _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2347_ _0253_ _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2278_ u_arbiter.i_wb_cpu_rdt\[15\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\]
+ u_cpu.cpu.genblk1.align.ctrl_misal _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2087__A1 _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3020__CLK net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3170__CLK net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2314__A2 u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2677__B _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[8\]_SI u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_cpu.rf_ram.RAM0_A[1] u_cpu.rf_ram.addr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xu_scanchain_local.scan_flop\[65\] u_scanchain_local.module_data_in\[64\] net145 u_arbiter.o_wb_cpu_adr\[27\]
+ net33 u_scanchain_local.module_data_in\[65\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2250__A1 _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1580_ u_cpu.cpu.immdec.imm19_12_20\[8\] _1027_ _1055_ u_cpu.cpu.immdec.imm24_20\[4\]
+ _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2201_ _0382_ _0383_ _0063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3181_ _0202_ net65 u_cpu.cpu.genblk3.csr.mcause3_0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2132_ u_arbiter.i_wb_cpu_dbus_dat\[3\] _0314_ _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2069__A1 _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2063_ _0270_ _0276_ _0031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3043__CLK net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2965_ _1260_ _1004_ _0282_ _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2241__A1 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2896_ _0561_ _0534_ _0960_ _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1916_ _1345_ u_cpu.rf_ram.i_wdata\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2792__A2 _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1847_ _1025_ _1288_ _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3193__CLK net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1778_ u_cpu.cpu.decode.opcode\[2\] _1031_ u_cpu.cpu.csr_d_sel _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_131_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3379_ u_scanchain_local.clk_out net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1807__A1 u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2535__A2 _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2299__A1 _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1897__I1 u_cpu.rf_ram.data\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3066__CLK net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2750_ _0859_ _0136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_fanout137_I net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1701_ u_arbiter.i_wb_cpu_dbus_adr\[19\] _1130_ _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2774__A2 _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2681_ _0414_ _0774_ _0814_ _0456_ _0817_ _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_12_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1632_ _1094_ _1102_ _1103_ u_arbiter.o_wb_cpu_adr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2526__A2 _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1563_ _1029_ _1037_ _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_28_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3164_ _0185_ net87 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3095_ _0120_ net111 u_arbiter.i_wb_cpu_dbus_adr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2115_ _0313_ _0315_ _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2046_ u_arbiter.i_wb_cpu_dbus_dat\[6\] _0262_ _0258_ _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_39_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2462__A1 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout27 net29 net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout16 net18 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout38 u_scanchain_local.clk net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout49 net50 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__2214__A1 u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2272__S _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2948_ u_cpu.cpu.genblk3.csr.mcause3_0\[2\] _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2879_ _0611_ _0619_ _0945_ _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2071__I _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2004__C _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2517__A2 _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2453__B2 _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2910__S _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2508__A2 _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[28\] u_arbiter.i_wb_cpu_rdt\[25\] net130 u_arbiter.i_wb_cpu_dbus_dat\[22\]
+ net16 u_arbiter.i_wb_cpu_rdt\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_37_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2156__I _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2802_ _0893_ _0154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_34_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2733_ _0850_ _0128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2664_ _0529_ _0797_ _0802_ _0412_ _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1615_ _1089_ _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2595_ _0459_ _0634_ _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1546_ u_cpu.cpu.bufreg.lsb\[1\] _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_8_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3216_ u_cpu.rf_ram_if.wdata1_r\[5\] net44 u_cpu.rf_ram_if.wdata1_r\[4\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3147_ _0169_ net117 u_cpu.cpu.ctrl.o_ibus_adr\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2683__A1 _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3078_ _0103_ net56 u_cpu.cpu.immdec.imm19_12_20\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2029_ _0246_ _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2435__A1 _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[17\]_SE net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2123__B1 _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2426__A1 _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2977__A2 _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3104__CLK net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[31\]_D u_arbiter.i_wb_cpu_rdt\[28\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2579__C _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2380_ _0494_ _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3001_ _0001_ net63 u_cpu.rf_ram_if.rdata0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1640__A2 _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[22\]_D u_arbiter.i_wb_cpu_rdt\[19\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_2716_ u_arbiter.i_wb_cpu_dbus_adr\[10\] u_arbiter.i_wb_cpu_dbus_adr\[11\] _0837_
+ _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2647_ _0766_ _0618_ _0698_ _0786_ _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2578_ _0562_ _0524_ _0569_ _0724_ _0549_ _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_43_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2656__A1 u_cpu.cpu.immdec.imm19_12_20\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2408__A1 _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1849__B _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2959__A2 _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1631__A2 _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[13\]_D u_arbiter.i_wb_cpu_rdt\[10\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2431__I1 u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2895__A1 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_cpu.rf_ram.RAM0_D[1] u_cpu.rf_ram.i_wdata\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1603__I u_cpu.cpu.genblk1.align.ctrl_misal vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2647__A1 _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xserv_0_157 io_oeb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1622__A2 _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1880_ _1271_ _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2501_ _0578_ _0649_ _0654_ _0634_ _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_68_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2432_ _0454_ _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2102__C _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2363_ _0473_ _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[40\]_CLK net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2294_ _0419_ _0462_ _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2638__A1 _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[55\]_CLK net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout32_I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2344__I _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2877__A1 _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2877__B2 _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2629__A1 _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[10\] u_arbiter.i_wb_cpu_rdt\[7\] net135 u_arbiter.i_wb_cpu_dbus_dat\[4\]
+ net21 u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__1915__I0 u_cpu.rf_ram_if.wdata0_r\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2981_ _1027_ _1014_ _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3200__D u_cpu.rf_ram_if.wdata0_r\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1932_ u_cpu.rf_ram_if.rdata1\[1\] _1354_ _1355_ _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1863_ _1239_ _1302_ _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1794_ _1028_ _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2020__A2 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2415_ _0564_ _0575_ _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2859__A1 u_cpu.cpu.ctrl.o_ibus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2346_ _0499_ _0504_ _0512_ _0079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2277_ _0249_ u_arbiter.i_wb_cpu_rdt\[14\] _0445_ _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_42_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2547__B1 _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2023__B _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_cpu.rf_ram.RAM0_A[0] u_cpu.rf_ram.addr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_58_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1589__A1 _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2786__B1 _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2250__A2 _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_scanchain_local.scan_flop\[58\] u_scanchain_local.module_data_in\[57\] net142 u_arbiter.o_wb_cpu_adr\[20\]
+ net27 u_scanchain_local.module_data_in\[58\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1761__A1 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2200_ u_arbiter.i_wb_cpu_rdt\[18\] _0380_ _0371_ u_arbiter.i_wb_cpu_dbus_dat\[18\]
+ _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2587__C _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3180_ _0201_ net67 u_cpu.cpu.genblk3.csr.mcause3_0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2159__I _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2131_ _0330_ _0046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2062_ u_cpu.raddr\[1\] _0273_ _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1998__I _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1816__A2 _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2108__B u_cpu.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2964_ _1248_ _0281_ _1003_ _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1915_ u_cpu.rf_ram_if.wdata0_r\[2\] u_cpu.rf_ram_if.wdata1_r\[2\] _1342_ _1345_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_120_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2241__A2 _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2895_ _0501_ _0603_ _0959_ _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2529__B1 _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1846_ _1269_ _1274_ _1277_ u_cpu.cpu.state.stage_two_req _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
X_1777_ u_arbiter.i_wb_cpu_dbus_we _1219_ u_cpu.cpu.immdec.imm24_20\[0\] _1221_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1752__A1 u_cpu.cpu.ctrl.o_ibus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[50\]_SE net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2329_ _0473_ _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_73_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2299__A2 _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2908__S _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[3\] u_arbiter.i_wb_cpu_rdt\[0\] net135 u_arbiter.i_wb_cpu_dbus_sel\[1\]
+ net22 u_arbiter.i_wb_cpu_rdt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_1_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1700_ _1155_ _1156_ _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2680_ _0254_ _0816_ _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1631_ u_arbiter.i_wb_cpu_dbus_adr\[5\] _1091_ _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1982__A1 u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1562_ _1040_ u_cpu.cpu.decode.op26 _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input4_I io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3163_ _0184_ net87 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2114_ _1317_ _0314_ _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3094_ _0119_ net107 u_arbiter.i_wb_cpu_dbus_adr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2045_ _1217_ _1276_ _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout28 net29 net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout17 net18 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__2462__A2 _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout39 u_arbiter.i_wb_cpu_dbus_dat\[1\] net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3160__CLK net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2214__A2 _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2947_ _0986_ _0989_ _0991_ _1051_ _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_fanout9_I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2878_ _0417_ _0495_ _0634_ _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__1973__A1 u_cpu.cpu.immdec.imm11_7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1829_ u_cpu.cpu.decode.opcode\[0\] _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2020__C _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2150__A1 u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2453__A2 _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2205__A2 _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1559__A4 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3033__CLK net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2692__A2 _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3183__CLK net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2801_ u_cpu.cpu.ctrl.o_ibus_adr\[9\] _0892_ _0887_ _1124_ _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2732_ u_arbiter.i_wb_cpu_dbus_adr\[17\] u_arbiter.i_wb_cpu_dbus_adr\[18\] _0849_
+ _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2663_ _0529_ _0800_ _0801_ _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1614_ _1088_ _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2594_ _0251_ u_arbiter.i_wb_cpu_rdt\[7\] _0739_ _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1545_ u_cpu.cpu.bufreg.lsb\[0\] _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3215_ u_cpu.rf_ram_if.wdata1_r\[4\] net43 u_cpu.rf_ram_if.wdata1_r\[3\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3146_ _0168_ net119 u_cpu.cpu.ctrl.o_ibus_adr\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout62_I net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3077_ _0102_ net55 u_cpu.cpu.immdec.imm19_12_20\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2347__I _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2028_ net2 _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3056__CLK net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2371__A1 _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2123__A1 u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2458__S _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2921__S _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2720__I _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[40\] u_scanchain_local.module_data_in\[39\] net138 u_arbiter.o_wb_cpu_adr\[2\]
+ net23 u_scanchain_local.module_data_in\[40\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_6_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3000_ _0000_ net63 u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2715_ _0840_ _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3079__CLK net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2646_ _0420_ _0519_ _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2577_ _0524_ _0425_ _0562_ _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2278__S u_cpu.cpu.genblk1.align.ctrl_misal vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3129_ _0151_ net107 u_cpu.cpu.ctrl.o_ibus_adr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2408__A2 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2026__B _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2592__A1 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2895__A2 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_cpu.rf_ram.RAM0_D[0] u_cpu.rf_ram.i_wdata\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2647__A2 _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xserv_0_158 io_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout112_I net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2500_ _0524_ _0579_ _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2431_ u_arbiter.i_wb_cpu_rdt\[21\] u_arbiter.i_wb_cpu_rdt\[5\] _0590_ _0591_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2362_ _0500_ _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2293_ _0250_ u_arbiter.i_wb_cpu_rdt\[8\] _0461_ _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_110_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[1\]_SE net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1861__A3 _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2810__A2 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout25_I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2629_ _0417_ _0617_ _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2877__A2 _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[14\]_SI u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2736__S _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2801__A2 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1614__I _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2980_ _1214_ _1014_ _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1931_ u_cpu.rf_ram_if.rtrig1 _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1862_ _1239_ _1302_ u_cpu.cpu.bne_or_bge _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1793_ _1035_ _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2414_ _0424_ _0543_ _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2859__A2 _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2345_ _1320_ _0505_ _0441_ _0511_ _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2276_ _0248_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[14\] _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_38_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2547__B2 _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2547__A1 _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2180__C1 _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_106_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2786__B2 u_cpu.cpu.ctrl.o_ibus_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2250__A3 _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[54\]_CLK net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2868__C _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1761__A2 u_cpu.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2130_ u_arbiter.i_wb_cpu_rdt\[1\] _0318_ _0329_ _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2884__B _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[69\]_CLK net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2061_ _0275_ _0030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2474__B1 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2108__C u_cpu.cpu.bufreg.lsb\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2226__B1 _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2963_ u_cpu.cpu.decode.co_ebreak _1246_ _1315_ _1245_ _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_37_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1914_ _1344_ u_cpu.rf_ram.i_wdata\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2777__A1 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2894_ _0429_ _0580_ _0593_ _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_33_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1845_ u_cpu.cpu.ctrl.pc_plus_offset_cy_r _1286_ _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2529__B2 _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1776_ u_arbiter.i_wb_cpu_dbus_we _1218_ _1219_ _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_144_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_fanout92_I net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2328_ _0484_ _0494_ _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2259_ u_arbiter.i_wb_cpu_rdt\[0\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\] _0427_
+ _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1807__A3 u_cpu.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2768__A1 _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2969__B _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2688__C _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1630_ _1100_ _1101_ _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1561_ u_cpu.cpu.decode.op21 _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_28_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3162_ _0183_ net82 u_cpu.cpu.genblk1.align.ctrl_misal vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2113_ _0258_ _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3093_ _0118_ net107 u_arbiter.i_wb_cpu_dbus_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2044_ u_arbiter.i_wb_cpu_dbus_dat\[5\] _0260_ _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_126_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1670__A1 u_arbiter.i_wb_cpu_dbus_adr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout29 net36 net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout18 net19 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_31_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2946_ _1033_ _1204_ u_cpu.cpu.genblk3.csr.mcause3_0\[2\] _1046_ _0988_ _0991_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_2877_ _0528_ _0441_ _0544_ _0545_ _0664_ _0703_ _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_50_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1973__A2 _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1828_ u_cpu.cpu.decode.co_mem_word _1028_ _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_117_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1759_ _1203_ _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1913__S _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2919__S _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout142_I net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2800_ _0875_ _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2731_ _1288_ _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_u_scanchain_local.scan_flop\[40\]_SE net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2601__B1 _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2662_ _0703_ _0578_ _0548_ _0797_ _0656_ _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
Xu_scanchain_local.output_buffers\[2\] u_scanchain_local.data_out_i u_scanchain_local.data_out
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2593_ _1080_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[7\] _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1613_ _1072_ u_cpu.cpu.state.ibus_cyc _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1707__A2 _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2904__A1 _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1544_ _1024_ u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_119_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3214_ u_cpu.rf_ram_if.wdata1_r\[3\] net41 u_cpu.rf_ram_if.wdata1_r\[2\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3145_ _0167_ net119 u_cpu.cpu.ctrl.o_ibus_adr\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1891__A1 _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout55_I net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3076_ _0101_ net56 u_cpu.cpu.immdec.imm19_12_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2027_ _0216_ _0245_ _0215_ u_arbiter.i_wb_cpu_dbus_sel\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2199__A2 _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2443__I0 u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2929_ _0980_ _0194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2371__A2 _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2123__A2 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[63\]_SE net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1937__A2 _0020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3000__CLK net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[33\] u_arbiter.i_wb_cpu_rdt\[30\] net144 u_arbiter.i_wb_cpu_dbus_dat\[27\]
+ net30 u_arbiter.i_wb_cpu_rdt\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__3150__CLK net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2822__B1 _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1625__A1 u_cpu.cpu.ctrl.o_ibus_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2183__I _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2714_ u_arbiter.i_wb_cpu_dbus_adr\[9\] u_arbiter.i_wb_cpu_dbus_adr\[10\] _0837_
+ _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2645_ _0545_ _0464_ _0467_ _0458_ _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2576_ u_arbiter.i_wb_cpu_rdt\[30\] u_arbiter.i_wb_cpu_rdt\[14\] _0590_ _0723_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3128_ _0150_ net107 u_cpu.cpu.ctrl.o_ibus_adr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3059_ _0084_ net66 u_cpu.cpu.csr_d_sel vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2813__B1 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3023__CLK net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2041__A1 _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3173__CLK net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1881__B _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1698__A4 _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1855__A1 _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xserv_0_159 io_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2804__B1 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2932__S _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2280__A1 _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2731__I _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout105_I net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2430_ _0589_ _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_68_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2361_ _0465_ _0495_ _0526_ _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_29_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2292_ _1078_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[8\] _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_2_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3214__D u_cpu.rf_ram_if.wdata1_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3046__CLK net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2271__A1 _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout18_I net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3196__CLK net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2023__A1 _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2641__I _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2326__A2 u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2628_ _0656_ _0557_ _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2559_ _0703_ _0557_ _0707_ _0664_ _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_82_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1921__S _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2037__B _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2262__A1 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3069__CLK net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1930_ _1353_ _0018_ _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1861_ _1258_ _1239_ _1302_ _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_35_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2005__A1 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2461__I _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1792_ u_cpu.cpu.bne_or_bge _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_66_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2413_ _0475_ _0482_ _0534_ _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2344_ _0510_ _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2275_ _0436_ _0438_ _0443_ _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_77_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2547__A2 _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2180__B1 _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2483__A1 _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2060_ _0255_ _0269_ _0273_ _0274_ _0275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__2474__A1 _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2474__B2 _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2962_ u_cpu.cpu.genblk3.csr.mie_mtie _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1913_ u_cpu.rf_ram_if.wdata0_r\[1\] u_cpu.rf_ram_if.wdata1_r\[1\] _1342_ _1344_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2405__B _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1985__B1 _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2893_ _0587_ _0954_ _0958_ _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1844_ _1285_ _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_129_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1775_ u_cpu.cpu.decode.opcode\[2\] u_cpu.cpu.decode.opcode\[0\] u_cpu.cpu.decode.opcode\[1\]
+ _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_98_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout85_I net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2327_ _0446_ _0493_ _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2258_ _0416_ _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2189_ _0345_ _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2465__A1 _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[1\]_D u_cpu.cpu.genblk3.csr.i_mtip vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2456__A1 _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xu_scanchain_local.scan_flop\[63\] u_scanchain_local.module_data_in\[62\] net145 u_arbiter.o_wb_cpu_adr\[25\]
+ net33 u_scanchain_local.module_data_in\[63\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1560_ u_cpu.cpu.decode.co_ebreak _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_67_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3161_ _0182_ net77 u_cpu.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2112_ _0312_ _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3092_ _0117_ net108 u_arbiter.i_wb_cpu_dbus_adr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2043_ u_arbiter.i_wb_cpu_dbus_dat\[4\] _0259_ _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout19 net20 net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__1670__A2 _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2945_ _0990_ _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2876_ _0940_ _0943_ _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1973__A3 _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1827_ u_cpu.cpu.genblk3.csr.o_new_irq u_cpu.cpu.state.genblk1.misalign_trap_sync_r
+ _1031_ _1268_ _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_11_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1758_ _1202_ _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1689_ _1149_ u_arbiter.o_wb_cpu_adr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2824__I _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[53\]_CLK net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[68\]_CLK net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1884__B _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2677__A1 _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[34\]_D u_arbiter.i_wb_cpu_rdt\[31\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2730_ _0848_ _0127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout135_I net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2601__B2 _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2661_ _0417_ _0776_ _0798_ _0771_ _0799_ _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_9_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1612_ _1075_ _1086_ _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2592_ _0592_ _0736_ _0737_ _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2365__B1 _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1543_ _1023_ _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3213_ u_cpu.rf_ram_if.wdata1_r\[2\] net40 u_cpu.rf_ram_if.wdata1_r\[1\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3144_ _0166_ net119 u_cpu.cpu.ctrl.o_ibus_adr\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3075_ _0100_ net61 u_cpu.cpu.immdec.imm7 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2026_ _1025_ _0216_ _0215_ u_arbiter.i_wb_cpu_dbus_sel\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout48_I net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[25\]_D u_arbiter.i_wb_cpu_rdt\[22\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2443__I1 u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2928_ u_arbiter.i_wb_cpu_rdt\[26\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[10\]
+ _0979_ _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2859_ u_cpu.cpu.ctrl.o_ibus_adr\[31\] _0876_ _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2659__A1 _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2755__S _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2554__I _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[16\]_D u_arbiter.i_wb_cpu_rdt\[13\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_scanchain_local.scan_flop\[26\] u_arbiter.i_wb_cpu_rdt\[23\] net129 u_arbiter.i_wb_cpu_dbus_dat\[20\]
+ net15 u_arbiter.i_wb_cpu_rdt\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_135_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2464__I _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2713_ _0839_ _0119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2644_ _0421_ _0578_ _0656_ _0556_ _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2575_ _0511_ _0715_ _0721_ _0498_ _0722_ _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_105_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2889__A1 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1543__I _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3127_ _0149_ net105 u_cpu.cpu.ctrl.o_ibus_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3058_ _0083_ net66 u_cpu.cpu.decode.co_mem_word vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2009_ u_cpu.cpu.ctrl.pc_plus_offset_cy_r _1286_ _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1919__S _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1718__I _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2041__A2 _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2280__A2 _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2360_ _0519_ _0525_ _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2291_ _0458_ _0459_ _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2099__A2 _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2271__A2 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2559__B1 _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2143__B _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1782__A1 _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2627_ _0622_ _0619_ _0767_ _0456_ _0768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA_u_scanchain_local.scan_flop\[53\]_SE net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2558_ u_arbiter.i_wb_cpu_rdt\[28\] u_arbiter.i_wb_cpu_rdt\[12\] _0589_ _0707_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_47_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2489_ _0644_ _0640_ _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2798__B1 _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2262__A2 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3140__CLK net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1828__A2 _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2789__B1 _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2742__I _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2253__A2 _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1860_ _1226_ _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2005__A2 _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1791_ _1066_ _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_7_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1764__A1 _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2412_ u_arbiter.i_wb_cpu_rdt\[20\] u_arbiter.i_wb_cpu_rdt\[4\] _1082_ _0573_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2189__I _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2343_ _0410_ _0509_ _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_96_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2274_ _0440_ _0441_ _0442_ _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_42_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2477__C1 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3013__CLK net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2229__C1 _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout30_I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3163__CLK net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1989_ _0215_ _0216_ _1037_ _1267_ _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_14_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2180__A1 u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1932__S _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2827__I _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2483__A2 _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_58_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1994__A1 _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1746__A1 _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3036__CLK net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2546__I0 u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2938__S _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3186__CLK net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2474__A2 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2226__A2 _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2961_ _1001_ _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1912_ _1343_ u_cpu.rf_ram.i_wdata\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1985__B2 _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2892_ _0587_ _0957_ _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1843_ _1219_ _1283_ _1284_ u_arbiter.i_wb_cpu_ibus_adr\[0\] _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__1737__A1 u_arbiter.i_wb_cpu_dbus_adr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1774_ u_cpu.cpu.immdec.imm11_7\[0\] _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_144_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2326_ _0250_ u_arbiter.i_wb_cpu_rdt\[15\] _0492_ _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout78_I net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2257_ _0422_ _0425_ _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2188_ _0373_ _0374_ _0059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2465__A2 _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1976__A1 u_cpu.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3059__CLK net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2528__I0 u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2456__A2 _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2208__A2 _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xu_scanchain_local.scan_flop\[56\] u_scanchain_local.module_data_in\[55\] net143 u_arbiter.o_wb_cpu_adr\[18\]
+ net29 u_scanchain_local.module_data_in\[56\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_32_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2392__A1 _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2668__S _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3160_ _0181_ net49 u_cpu.cpu.immdec.imm11_7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3091_ _0116_ net108 u_arbiter.i_wb_cpu_dbus_adr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2467__I _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2111_ _0256_ _0311_ _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2042_ u_arbiter.i_wb_cpu_dbus_dat\[3\] u_arbiter.i_wb_cpu_dbus_dat\[2\] u_arbiter.i_wb_cpu_dbus_dat\[0\]
+ net39 _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_48_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2447__A2 _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2944_ _0987_ u_cpu.cpu.genblk3.csr.mcause3_0\[0\] _0989_ _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2875_ _0695_ _0511_ _0942_ _0489_ _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3201__CLK net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1826_ u_cpu.cpu.genblk3.csr.o_new_irq u_cpu.cpu.state.init_done _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__2383__A1 _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1757_ _1200_ _1201_ _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_117_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1688_ u_arbiter.i_wb_cpu_dbus_adr\[16\] _1148_ _1074_ _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2135__A1 u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2930__I0 u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2309_ _0456_ _0469_ _0474_ _0475_ _0477_ _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__2377__I _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1716__A4 _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2921__I0 u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2677__A2 _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_scanchain_local.scan_flop\[1\] u_cpu.cpu.genblk3.csr.i_mtip net139 u_arbiter.o_wb_cpu_we
+ net25 u_arbiter.i_wb_cpu_ack vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_92_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1652__A3 _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2601__A2 _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout128_I net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2660_ _0507_ _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_12_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1611_ _1083_ _1084_ _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2591_ _0621_ _0501_ _0534_ _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2365__B2 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2365__A1 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1542_ _1020_ _1021_ _1022_ _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_3212_ u_cpu.rf_ram_if.wdata1_r\[1\] net40 u_cpu.rf_ram_if.wdata1_r\[0\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2912__I0 u_arbiter.i_wb_cpu_rdt\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input2_I io_in[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3143_ _0165_ net119 u_cpu.cpu.ctrl.o_ibus_adr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3074_ _0099_ net73 u_cpu.cpu.immdec.imm30_25\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2025_ _1026_ _0245_ _0215_ u_arbiter.i_wb_cpu_dbus_sel\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_u_scanchain_local.scan_flop\[4\]_SE net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2927_ _0252_ _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2858_ _0923_ _0926_ _0927_ _1243_ _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_102_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2789_ u_cpu.cpu.ctrl.o_ibus_adr\[4\] _0885_ _0880_ _1100_ _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2356__A1 _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1809_ _1250_ _1251_ _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1954__I1 _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2659__A2 _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1634__A3 _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[19\] u_arbiter.i_wb_cpu_rdt\[16\] net127 u_arbiter.i_wb_cpu_dbus_dat\[13\]
+ net13 u_arbiter.i_wb_cpu_rdt\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_2_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1570__A2 _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2822__A2 _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2712_ u_arbiter.i_wb_cpu_dbus_adr\[8\] u_arbiter.i_wb_cpu_dbus_adr\[9\] _0837_ _0839_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2586__A1 _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2643_ _0548_ _0782_ _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2574_ u_cpu.cpu.immdec.imm30_25\[4\] _0685_ _0711_ u_cpu.cpu.immdec.imm30_25\[5\]
+ _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_82_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2889__A2 _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1824__I _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3126_ _0148_ net105 u_cpu.cpu.ctrl.o_ibus_adr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout60_I net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2510__A1 _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[67\]_CLK net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3057_ _0082_ net66 u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2813__A2 _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2008_ _0226_ _0232_ _0233_ _0014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2577__A1 _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2604__B _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1935__S _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2501__A1 _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2804__A2 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2568__A1 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2290_ u_arbiter.i_wb_cpu_rdt\[13\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[13\]
+ _1078_ _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2559__A1 _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1819__I _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2559__B2 _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2626_ _0438_ _0465_ _0766_ _0619_ _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__1782__A2 _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3092__CLK net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2557_ _0703_ _0484_ _0544_ _0553_ _0705_ _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_88_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2488_ u_cpu.cpu.immdec.imm24_20\[1\] _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_29_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3109_ _0134_ net120 u_arbiter.i_wb_cpu_dbus_adr\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2509__B _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2789__A1 u_cpu.cpu.ctrl.o_ibus_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1639__I _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1790_ _1233_ _0013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout110_I net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2411_ _1029_ _0515_ _0572_ _0084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2342_ _0506_ _0507_ _0508_ _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2273_ u_arbiter.i_wb_cpu_rdt\[2\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[2\] _0427_
+ _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2477__B1 _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2477__C2 _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2229__B1 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout23_I net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[20\]_SE net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1988_ _1026_ _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2601__C _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2609_ _1232_ _0753_ _0513_ _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2180__A2 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_58_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2546__I1 u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2960_ u_cpu.cpu.genblk3.csr.mstatus_mie u_cpu.cpu.genblk3.csr.mstatus_mpie _1000_
+ _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_u_scanchain_local.scan_flop\[43\]_SE net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2891_ _0457_ _0603_ _0549_ _0517_ _0956_ _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1911_ u_cpu.rf_ram_if.wdata0_r\[0\] u_cpu.rf_ram_if.wdata1_r\[0\] _1342_ _1343_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1842_ _1271_ u_cpu.cpu.decode.opcode\[1\] _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_129_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1737__A2 _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1773_ u_cpu.cpu.bufreg2.i_cnt_done _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2325_ _1078_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\] _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3130__CLK net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2256_ _0424_ _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2187_ u_arbiter.i_wb_cpu_rdt\[14\] _0364_ _0371_ u_arbiter.i_wb_cpu_dbus_dat\[14\]
+ _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_129_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2870__B1 _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1976__A2 _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2998__CLK net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1728__A2 _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2528__I1 u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2689__B1 _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[66\]_SE net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1719__A2 _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[49\] u_scanchain_local.module_data_in\[48\] net141 u_arbiter.o_wb_cpu_adr\[11\]
+ net27 u_scanchain_local.module_data_in\[49\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_67_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2392__A2 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3153__CLK net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3090_ _0115_ net106 u_arbiter.i_wb_cpu_dbus_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2110_ _1231_ _0309_ _0310_ _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2041_ _0256_ _0257_ _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_78_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2943_ _0988_ _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_16_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2874_ _1386_ _0930_ _0941_ _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1825_ _1025_ _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1756_ u_cpu.rf_ram_if.rcnt\[0\] _1021_ _1022_ u_cpu.rf_ram_if.wen0_r _1201_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_144_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2383__A2 _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1687_ _1147_ _1145_ _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_fanout90_I net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2308_ _0476_ _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2686__A3 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2239_ _0406_ _0394_ _0354_ _1302_ _0408_ _0076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3026__CLK net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1938__S _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2342__B _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2921__I1 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1885__A1 _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2834__B1 _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1647__I _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1610_ _1083_ _1084_ _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2590_ _0419_ _0421_ _0425_ _0449_ _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__2365__A2 _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1541_ u_cpu.rf_ram_if.rcnt\[1\] _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_10_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3211_ _0214_ net64 u_cpu.rf_ram_if.rcnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3142_ _0164_ net115 u_cpu.cpu.ctrl.o_ibus_adr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3073_ _0098_ net75 u_cpu.cpu.immdec.imm30_25\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2825__B1 _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_cpu.rf_ram.RAM0_CLK net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2024_ _1235_ _1025_ _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3049__CLK net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2926_ _0978_ _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3199__CLK net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2053__A1 _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1800__A1 _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2857_ _0923_ _1307_ _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1808_ _1217_ u_cpu.cpu.genblk3.csr.mcause31 _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2788_ _0876_ _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1739_ u_cpu.cpu.ctrl.o_ibus_adr\[27\] _1181_ _1182_ _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_46_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2388__I _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2108__A2 u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1867__A1 _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2816__B1 _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2337__B _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2292__A1 _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2044__A1 u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2595__A2 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2072__B _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.output_buffers\[3\]_I net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2658__I0 u_arbiter.i_wb_cpu_rdt\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2283__A1 _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2035__A1 _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout140_I net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2711_ _0838_ _0118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2642_ u_arbiter.i_wb_cpu_rdt\[16\] u_arbiter.i_wb_cpu_rdt\[0\] _0589_ _0782_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_127_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2573_ _0654_ _0716_ _0720_ _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1849__A1 u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3125_ _0147_ net105 u_cpu.cpu.ctrl.o_ibus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout53_I net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3056_ _0081_ net60 u_cpu.cpu.branch_op vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2007_ _1279_ _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_24_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2909_ _0969_ _0185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2501__A2 _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2265__A1 _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2514__C _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_scanchain_local.scan_flop\[31\] u_arbiter.i_wb_cpu_rdt\[28\] net131 u_arbiter.i_wb_cpu_dbus_dat\[25\]
+ net17 u_arbiter.i_wb_cpu_rdt\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_2_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2559__A2 _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2625_ _0552_ _0483_ _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1782__A3 _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2556_ _0626_ _0704_ _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2487_ _0639_ _0642_ _0643_ _0586_ _0089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_130_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3108_ _0133_ net119 u_arbiter.i_wb_cpu_dbus_adr\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3039_ _0064_ net99 u_arbiter.i_wb_cpu_dbus_dat\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2798__A2 _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2486__A1 u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2238__A1 u_arbiter.i_wb_cpu_rdt\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2789__A2 _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[66\]_CLK net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1655__I _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout103_I net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2410_ _0568_ _0571_ _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2174__B1 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2687__S _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2341_ _0453_ _0432_ _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_96_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2272_ u_arbiter.i_wb_cpu_rdt\[4\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[4\] _0427_
+ _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2477__B2 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2477__A1 _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2229__A1 u_arbiter.i_wb_cpu_rdt\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[19\]_CLK net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2435__B _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout16_I net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1987_ _1236_ _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2401__A1 _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2608_ _1222_ _1292_ _0752_ _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2539_ _0254_ _0684_ _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2468__A1 _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_106_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[4\]_D u_arbiter.i_wb_cpu_rdt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2459__A1 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2890_ _0799_ _0951_ _0955_ _0415_ _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_31_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1910_ _1341_ _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__2631__A1 _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1841_ _1264_ u_arbiter.i_wb_cpu_dbus_we _1039_ _1049_ _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1772_ u_cpu.rf_ram_if.rdata1\[0\] _1214_ _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2324_ _0470_ _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2255_ u_arbiter.i_wb_cpu_rdt\[12\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[12\]
+ _0423_ _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2186_ u_arbiter.i_wb_cpu_dbus_dat\[15\] _0358_ _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2870__A1 _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2870__B2 _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2622__A1 u_cpu.cpu.csr_imm vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2689__A1 u_cpu.cpu.immdec.imm31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2310__B1 _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2854__I _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2861__A1 _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[46\]_D u_scanchain_local.module_data_in\[45\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2040_ _1268_ _1273_ _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_u_scanchain_local.scan_flop\[10\]_SE net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2604__A1 _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2942_ _0277_ _1052_ _1254_ _1247_ _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_31_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2873_ u_cpu.cpu.immdec.imm11_7\[1\] _0930_ _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_11_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1824_ _1265_ _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1755_ u_cpu.rf_ram_if.wen1_r u_cpu.rf_ram_if.genblk1.wtrig0_r _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1686_ u_cpu.cpu.ctrl.o_ibus_adr\[16\] _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_fanout83_I net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2540__B1 _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2307_ _0410_ _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2238_ u_arbiter.i_wb_cpu_rdt\[31\] _0267_ _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1646__A2 _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2169_ _0345_ _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[28\]_D u_arbiter.i_wb_cpu_rdt\[25\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1954__S u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[33\]_SE net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2382__I0 u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_u_scanchain_local.scan_flop\[19\]_D u_arbiter.i_wb_cpu_rdt\[16\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1928__I u_cpu.rf_ram.regzero vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_scanchain_local.scan_flop\[61\] u_scanchain_local.module_data_in\[60\] net145 u_arbiter.o_wb_cpu_adr\[23\]
+ net33 u_scanchain_local.module_data_in\[61\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_139_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3120__CLK net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1540_ u_cpu.rf_ram_if.rcnt\[2\] _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_5_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2759__I u_arbiter.i_wb_cpu_dbus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3210_ u_cpu.rf_ram_if.rtrig0 net52 u_cpu.rf_ram_if.rtrig1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3141_ _0163_ net114 u_cpu.cpu.ctrl.o_ibus_adr\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2695__S _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3072_ _0097_ net61 u_cpu.cpu.immdec.imm30_25\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2023_ _1234_ _0244_ _0219_ u_cpu.cpu.o_wen0 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_78_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2925_ u_arbiter.i_wb_cpu_rdt\[25\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[9\]
+ _0973_ _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2053__A2 _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1800__A2 _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2856_ u_cpu.cpu.ctrl.i_jump _1296_ _0925_ _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_15_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1807_ u_cpu.cpu.mem_bytecnt\[1\] u_cpu.cpu.state.o_cnt\[2\] u_cpu.cpu.mem_bytecnt\[0\]
+ _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_2787_ _0884_ _0148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_89_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[56\]_SE net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1738_ _1174_ _1186_ _1187_ u_arbiter.o_wb_cpu_adr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1669_ _1133_ _1129_ _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_59_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2513__B1 _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2292__A2 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3143__CLK net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1858__A2 _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2658__I1 u_arbiter.i_wb_cpu_rdt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2035__A2 u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2710_ u_arbiter.i_wb_cpu_dbus_adr\[7\] u_arbiter.i_wb_cpu_dbus_adr\[8\] _0837_ _0838_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2641_ _0757_ _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2572_ _0717_ _0719_ _0620_ _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_141_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3016__CLK net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3124_ _0146_ net81 u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3055_ _0080_ net73 u_arbiter.i_wb_cpu_dbus_we vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3166__CLK net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2006_ _0228_ _0231_ _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2274__A2 _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout46_I net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1568__I u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2026__A2 _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2908_ u_arbiter.i_wb_cpu_rdt\[17\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\]
+ _0967_ _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2839_ _0878_ _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2265__A2 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3039__CLK net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2576__I0 u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[24\] u_arbiter.i_wb_cpu_rdt\[21\] net128 u_arbiter.i_wb_cpu_dbus_dat\[18\]
+ net13 u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_29_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3189__CLK net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2624_ u_cpu.cpu.csr_imm _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_138_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2555_ _0605_ _0464_ _0627_ _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2486_ u_cpu.cpu.immdec.imm24_20\[0\] _0642_ _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3107_ _0132_ net115 u_arbiter.i_wb_cpu_dbus_adr\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3038_ _0063_ net99 u_arbiter.i_wb_cpu_dbus_dat\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2558__I0 u_arbiter.i_wb_cpu_rdt\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1962__S _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2486__A2 _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2238__A2 _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1749__A1 _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2410__A2 _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2174__A1 u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2340_ _0428_ _0454_ _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_81_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2271_ _1079_ _0337_ _0439_ _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2721__I0 u_arbiter.i_wb_cpu_dbus_adr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2477__A2 _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2229__A2 _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2435__C _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1986_ _1058_ net8 _1387_ u_cpu.rf_ram.addr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__2401__A2 _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2607_ _1310_ _0222_ _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2538_ _0681_ _0686_ _0689_ _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2469_ _0552_ _0463_ _0459_ _0458_ _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_69_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2626__B _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1691__A3 _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2640__A2 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2631__A2 _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1840_ _1281_ _1247_ _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1771_ _1210_ _1213_ u_cpu.rf_ram.regzero _1214_ _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__2395__A1 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2323_ _0413_ _0488_ _0490_ _0078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2254_ _0416_ _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2185_ _0370_ _0372_ _0058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_u_scanchain_local.scan_flop\[7\]_SE net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1673__A3 _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2870__A2 _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2622__A2 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1969_ u_cpu.raddr\[1\] _1378_ _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_135_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2689__A2 _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[50\]_CLK net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2310__B2 _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[65\]_CLK net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2861__A2 _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_u_cpu.rf_ram.RAM0_WEN[7] net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2613__A2 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[18\]_CLK net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2852__A2 _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2941_ _1045_ _0986_ _1051_ _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2604__A2 _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2872_ _0587_ _0939_ _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1823_ _1264_ _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1754_ _1075_ _1198_ _1199_ u_arbiter.o_wb_cpu_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1685_ _1122_ _1143_ _1145_ _1146_ u_arbiter.o_wb_cpu_adr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_144_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_fanout76_I net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2306_ _0442_ _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2237_ _0404_ _0394_ _0354_ _0406_ _0407_ _0075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_39_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2168_ _0359_ _0360_ _0053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2099_ u_cpu.cpu.alu.cmp_r _1307_ _1300_ _0298_ _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_59_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2906__I0 u_arbiter.i_wb_cpu_rdt\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3072__CLK net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2382__I1 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2531__A1 _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2834__A2 _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2598__A1 _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[54\] u_scanchain_local.module_data_in\[53\] net132 u_arbiter.o_wb_cpu_adr\[16\]
+ net18 u_scanchain_local.module_data_in\[54\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_138_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2770__A1 u_arbiter.i_wb_cpu_dbus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3140_ _0162_ net99 u_cpu.cpu.ctrl.o_ibus_adr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2522__A1 _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2775__I _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3071_ _0096_ net75 u_cpu.cpu.immdec.imm30_25\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2825__A2 _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2022_ u_cpu.cpu.immdec.imm11_7\[4\] _0241_ _0242_ _0243_ _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_91_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2589__A1 _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2924_ _0977_ _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2855_ u_cpu.cpu.ctrl.i_jump _0924_ _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1806_ _1244_ _1245_ _1247_ _1248_ _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_89_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2786_ u_cpu.cpu.ctrl.o_ibus_adr\[3\] _0877_ _0880_ u_cpu.cpu.ctrl.o_ibus_adr\[4\]
+ _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_116_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1737_ u_arbiter.i_wb_cpu_dbus_adr\[27\] _1172_ _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3095__CLK net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1668_ u_cpu.cpu.ctrl.o_ibus_adr\[12\] _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1599_ _1071_ _1075_ _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2513__A1 _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2513__B2 _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2816__A2 _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2634__B _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1555__A2 _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2504__A1 _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2640_ _0765_ _0756_ _0779_ _0780_ _0105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_139_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2571_ _0624_ _0718_ _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_5_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3123_ _0145_ net81 u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3054_ _0079_ net73 u_cpu.cpu.decode.opcode\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2005_ _1310_ _1224_ _0230_ _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_64_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2274__A3 _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[23\]_SE net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2907_ _0968_ _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2982__A1 _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2838_ _0914_ _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2769_ _1267_ _0870_ _0871_ _0143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[30\]_SI u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3110__CLK net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2273__I0 u_arbiter.i_wb_cpu_rdt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1695__S _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1776__A2 _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2973__A1 _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2576__I1 u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[17\] u_arbiter.i_wb_cpu_rdt\[14\] net128 u_arbiter.i_wb_cpu_dbus_dat\[11\]
+ net14 u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_42_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[46\]_SE net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2964__A1 _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2623_ _0763_ _0756_ _0764_ _0572_ _0104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2554_ _0417_ _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2485_ _0641_ _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3133__CLK net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3106_ _0131_ net114 u_arbiter.i_wb_cpu_dbus_adr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3037_ _0062_ net89 u_arbiter.i_wb_cpu_dbus_dat\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2255__I0 u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2558__I1 u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[69\]_SE net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2891__B1 _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1997__A2 _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2246__I0 u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3006__CLK net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2946__A1 _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2113__I _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2174__A2 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3156__CLK net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2270_ _0423_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[3\] _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1685__A1 _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2882__B1 _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1985_ _1059_ _1380_ _1385_ _1389_ u_cpu.rf_ram.addr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_53_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2606_ _0749_ _0750_ _0751_ _0219_ _0100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2537_ u_cpu.cpu.immdec.imm30_25\[0\] _0688_ _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2468_ _0593_ _0623_ _0625_ _0618_ _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_25_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2712__I1 u_arbiter.i_wb_cpu_dbus_adr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2399_ _0521_ _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1676__A1 u_arbiter.i_wb_cpu_dbus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2626__C _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_58_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_58_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3179__CLK net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1770_ u_cpu.rf_ram_if.rtrig1 _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_144_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2778__I _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2552__C1 _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2322_ _0222_ _0489_ _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2253_ _0419_ _0421_ _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2184_ u_arbiter.i_wb_cpu_rdt\[13\] _0364_ _0371_ u_arbiter.i_wb_cpu_dbus_dat\[13\]
+ _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2458__I0 u_arbiter.i_wb_cpu_rdt\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2462__B _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1968_ u_cpu.raddr\[0\] _1376_ _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1899_ u_cpu.rf_ram.rdata\[3\] u_cpu.rf_ram.data\[3\] _1333_ _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1649__A1 _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2310__A2 _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_cpu.rf_ram.RAM0_WEN[6] net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2074__A1 _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1888__A1 _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2837__B1 _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2940_ u_cpu.cpu.genblk3.csr.mcause3_0\[1\] _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_16_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2871_ _0934_ _0937_ _0938_ _0598_ _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1822_ _1031_ _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1753_ u_arbiter.i_wb_cpu_dbus_adr\[31\] _1074_ _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1684_ u_arbiter.i_wb_cpu_dbus_adr\[15\] _1130_ _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1591__A3 _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2540__A2 _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2305_ _0473_ _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2828__B1 _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2236_ u_arbiter.i_wb_cpu_rdt\[30\] _0267_ _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout69_I net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2167_ u_arbiter.i_wb_cpu_rdt\[8\] _0339_ _0348_ u_arbiter.i_wb_cpu_dbus_dat\[8\]
+ _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_54_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2098_ _1229_ _0301_ _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2359__A2 _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2412__S _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2211__I _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3217__CLK net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2531__A2 _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2367__B _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2047__A1 _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[47\] u_scanchain_local.module_data_in\[46\] net146 u_arbiter.o_wb_cpu_adr\[9\]
+ net27 u_scanchain_local.module_data_in\[47\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__2770__A2 _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3070_ _0095_ net75 u_cpu.cpu.immdec.imm30_25\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_u_scanchain_local.input_buf_clk_I net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2021_ _0237_ _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2791__I _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2038__A1 _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2923_ u_arbiter.i_wb_cpu_rdt\[24\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[8\]
+ _0973_ _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2854_ _1327_ _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2785_ _0883_ _0147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1805_ u_cpu.cpu.decode.op26 _1043_ _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1736_ u_cpu.cpu.ctrl.o_ibus_adr\[27\] _1185_ _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_102_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[64\]_CLK net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1667_ _1093_ _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2761__A2 _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1598_ _1074_ _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2513__A2 _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2219_ u_arbiter.i_wb_cpu_rdt\[24\] _0321_ _0352_ u_arbiter.i_wb_cpu_dbus_dat\[25\]
+ _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_45_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3199_ u_cpu.rf_ram_if.wdata0_r\[1\] net40 u_cpu.rf_ram_if.wdata0_r\[0\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[17\]_CLK net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2268__A1 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2116__I _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2440__A1 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout119_I net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2570_ _0618_ _0623_ _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3122_ _0015_ net80 u_cpu.cpu.ctrl.pc_plus_4_cy_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3053_ _0078_ net73 u_cpu.cpu.decode.opcode\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2004_ _0229_ _1284_ _1307_ _1265_ _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_91_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2906_ u_arbiter.i_wb_cpu_rdt\[16\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\]
+ _0967_ _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_17_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2837_ u_cpu.cpu.ctrl.o_ibus_adr\[24\] _0913_ _0908_ u_cpu.cpu.ctrl.o_ibus_adr\[25\]
+ _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2768_ _1026_ _0870_ _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1719_ u_arbiter.i_wb_cpu_dbus_adr\[23\] _1172_ _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2699_ u_arbiter.i_wb_cpu_dbus_adr\[2\] u_arbiter.i_wb_cpu_dbus_adr\[3\] _0831_ _0832_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2498__A1 _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2645__B _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2670__A1 _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3085__CLK net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2661__A1 _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2413__A1 _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2964__A2 _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2622_ u_cpu.cpu.csr_imm _0505_ _0757_ _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2177__B1 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2553_ _0701_ _0702_ _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2484_ _0476_ _0640_ _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3105_ _0130_ net114 u_arbiter.i_wb_cpu_dbus_adr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3036_ _0061_ net93 u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout51_I net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_cpu.rf_ram.RAM0_GWEN _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2652__A1 _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2404__A1 _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1595__I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2891__A1 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2891__B2 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2643__A1 _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2946__A2 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[7\]_D u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[13\]_SE net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2882__A1 u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1984_ u_cpu.cpu.immdec.imm11_7\[4\] _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA_u_scanchain_local.out_flop_CLKN net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3100__CLK net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2605_ u_cpu.cpu.immdec.imm7 _0542_ _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_fanout99_I net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2536_ _0254_ _0687_ _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2467_ _0624_ _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2398_ _0509_ _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1676__A2 _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2873__A1 u_cpu.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2625__A1 _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3019_ _0044_ net69 u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XPHY_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_106_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[36\]_SE net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3192__D _0020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout150 net151 net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__2864__A1 u_cpu.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2092__A2 _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout101_I net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2552__B1 _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2552__C2 _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2321_ _0411_ _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2252_ _0420_ _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2183_ _0322_ _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2607__A1 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2458__I1 u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1830__A2 _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout14_I net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1967_ _1377_ u_cpu.rf_ram.addr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_u_scanchain_local.scan_flop\[59\]_SE net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1898_ _1335_ _0019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1873__I u_cpu.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2519_ _0668_ _0671_ _0093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_cpu.rf_ram.RAM0_WEN[5] net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3146__CLK net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2653__B _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2074__A2 _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1585__A1 u_cpu.cpu.immdec.imm19_12_20\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2782__B1 _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2065__A2 _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout149_I net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2870_ _0528_ _0487_ _0664_ _0695_ _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1812__A2 _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1821_ _1261_ _1263_ u_cpu.cpu.o_wdata1 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1752_ u_cpu.cpu.ctrl.o_ibus_adr\[31\] _1195_ _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1576__A1 _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1683_ u_cpu.cpu.ctrl.o_ibus_adr\[13\] u_cpu.cpu.ctrl.o_ibus_adr\[12\] _1129_ _1144_
+ _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2304_ _0448_ _0471_ _0472_ _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2235_ u_arbiter.i_wb_cpu_dbus_dat\[31\] _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2166_ u_arbiter.i_wb_cpu_dbus_dat\[9\] _0358_ _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2029__I _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2097_ _1239_ _1302_ _0300_ _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_94_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2999_ _0012_ net51 u_cpu.rf_ram_if.rdata1\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xu_cpu.rf_ram.RAM0 u_cpu.rf_ram.RAM0/A[0] u_cpu.rf_ram.RAM0/A[1] u_cpu.rf_ram.RAM0/A[2]
+ u_cpu.rf_ram.RAM0/A[3] u_cpu.rf_ram.RAM0/A[4] u_cpu.rf_ram.RAM0/A[5] u_cpu.rf_ram.RAM0/A[6]
+ u_cpu.rf_ram.RAM0/A[7] u_cpu.rf_ram.RAM0/CEN u_cpu.rf_ram.RAM0/CLK u_cpu.rf_ram.RAM0/D[0]
+ u_cpu.rf_ram.RAM0/D[1] u_cpu.rf_ram.RAM0/D[2] u_cpu.rf_ram.RAM0/D[3] u_cpu.rf_ram.RAM0/D[4]
+ u_cpu.rf_ram.RAM0/D[5] u_cpu.rf_ram.RAM0/D[6] u_cpu.rf_ram.RAM0/D[7] u_cpu.rf_ram.RAM0/GWEN
+ u_cpu.rf_ram.RAM0/Q[0] u_cpu.rf_ram.RAM0/Q[1] u_cpu.rf_ram.RAM0/Q[2] u_cpu.rf_ram.RAM0/Q[3]
+ u_cpu.rf_ram.RAM0/Q[4] u_cpu.rf_ram.RAM0/Q[5] u_cpu.rf_ram.RAM0/Q[6] u_cpu.rf_ram.RAM0/Q[7]
+ u_cpu.rf_ram.RAM0/WEN[0] u_cpu.rf_ram.RAM0/WEN[1] u_cpu.rf_ram.RAM0/WEN[2] u_cpu.rf_ram.RAM0/WEN[3]
+ u_cpu.rf_ram.RAM0/WEN[4] u_cpu.rf_ram.RAM0/WEN[5] u_cpu.rf_ram.RAM0/WEN[6] u_cpu.rf_ram.RAM0/WEN[7]
+ vdd vss gf180mcu_fd_ip_sram__sram256x8m8wm1
XFILLER_134_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2020_ _1321_ _1204_ _1328_ _1310_ _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_78_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2286__A2 _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2038__A2 _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2922_ _0976_ _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2853_ _1052_ _0922_ _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_141_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2784_ _1084_ _0877_ _0880_ u_cpu.cpu.ctrl.o_ibus_adr\[3\] _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_15_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1804_ _1246_ u_cpu.cpu.state.o_cnt\[2\] u_cpu.cpu.mem_bytecnt\[0\] _1247_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_1735_ _1181_ _1182_ _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2312__I _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1666_ _1111_ _1127_ _1129_ _1131_ u_arbiter.o_wb_cpu_adr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1597_ _1073_ _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_131_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout81_I net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2218_ u_arbiter.i_wb_cpu_dbus_dat\[24\] _0394_ _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2277__A2 u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3198_ _0210_ net81 u_cpu.cpu.state.ibus_cyc vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2149_ _0345_ _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1598__I _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2512__I0 u_arbiter.i_wb_cpu_rdt\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2268__A2 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1779__A1 u_cpu.cpu.bufreg2.i_cnt_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1971__I _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3121_ _0016_ net80 u_cpu.cpu.ctrl.pc_plus_offset_cy_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3052_ _0077_ net73 u_cpu.cpu.decode.opcode\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2003_ _1321_ _0222_ _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_1_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2307__I _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3207__CLK net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2905_ _0252_ _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_32_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2836_ _0875_ _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2767_ _1279_ _0257_ _0869_ _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1718_ _1090_ _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2698_ _0830_ _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1649_ _1111_ _1114_ _1115_ _1117_ u_arbiter.o_wb_cpu_adr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_28_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2498__A2 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2217__I _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_109_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1791__I _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2489__A2 _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2110__A1 _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[63\]_CLK net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2661__A2 _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2413__A2 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout131_I net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2177__A1 u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2621_ u_cpu.cpu.immdec.imm19_12_20\[3\] _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_103_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2552_ u_cpu.cpu.immdec.imm30_25\[2\] _0688_ _0690_ u_cpu.cpu.immdec.imm30_25\[3\]
+ _0696_ _0588_ _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_142_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2483_ _0297_ _1209_ _1034_ _1232_ _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA_u_scanchain_local.scan_flop\[16\]_CLK net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3104_ _0129_ net114 u_arbiter.i_wb_cpu_dbus_adr\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3035_ _0060_ net89 u_arbiter.i_wb_cpu_dbus_dat\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2101__A1 _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout44_I net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2404__A2 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2819_ _0903_ _0161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_30_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2701__S _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2340__A1 _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2891__A2 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2643__A2 _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2391__B _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[22\] u_arbiter.i_wb_cpu_rdt\[19\] net127 u_arbiter.i_wb_cpu_dbus_dat\[16\]
+ net14 u_arbiter.i_wb_cpu_rdt\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_46_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3052__CLK net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1685__A3 _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2882__A2 _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1897__S _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1983_ _1056_ _1380_ _1388_ u_cpu.rf_ram.addr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_2604_ _0218_ _0732_ _0638_ _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2570__A1 _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2535_ _0297_ _0682_ _0218_ _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2466_ _0414_ _0523_ _0424_ _0518_ _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_87_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2322__A1 _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2397_ _0541_ _0515_ _0560_ _0082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2873__A2 _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2625__A2 _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3018_ _0043_ net79 u_cpu.cpu.bufreg2.i_cnt_done vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_58_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2431__S _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2936__I0 u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3075__CLK net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2561__A1 _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout140 net150 net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__2313__A1 _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout151 net4 net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__2386__B _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2864__A2 _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2616__A2 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2320_ _0456_ _0485_ _0474_ _0487_ _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2251_ u_arbiter.i_wb_cpu_rdt\[8\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[8\] _1079_
+ _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2304__A1 _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2182_ u_arbiter.i_wb_cpu_dbus_dat\[14\] _0358_ _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2607__A2 _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1966_ u_cpu.raddr\[0\] _1376_ _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__3098__CLK net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2251__S _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1897_ u_cpu.rf_ram.rdata\[2\] u_cpu.rf_ram.data\[2\] _1333_ _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[9\]_CLK net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2543__A1 _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2518_ u_cpu.cpu.immdec.imm24_20\[4\] _0641_ _0665_ _0588_ _0670_ _0671_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_97_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2449_ _0453_ _0454_ _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_cpu.rf_ram.RAM0_WEN[4] net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2782__A1 u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1585__A2 _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1820_ _1071_ _1262_ _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1751_ _1194_ _1196_ _1197_ u_arbiter.o_wb_cpu_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2773__A1 _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1682_ u_cpu.cpu.ctrl.o_ibus_adr\[15\] u_cpu.cpu.ctrl.o_ibus_adr\[14\] _1144_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_99_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2525__A1 _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2303_ _0429_ _0454_ _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2828__A2 _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2234_ _0403_ _0394_ _0354_ _0404_ _0405_ _0074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2165_ _0346_ _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2096_ _1238_ _1226_ _0299_ _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[26\]_SE net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2998_ _0011_ net51 u_cpu.rf_ram_if.rdata1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1949_ _1210_ _1213_ u_cpu.rf_ram.regzero _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_31_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2648__C _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3113__CLK net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1794__I _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[49\]_SE net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2921_ u_arbiter.i_wb_cpu_rdt\[23\] u_cpu.cpu.genblk1.align.ibus_rdt_concat\[7\]
+ _0973_ _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_44_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1797__A2 u_cpu.cpu.csr_imm vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2852_ _1040_ _1049_ _1042_ _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_102_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2783_ _0882_ _0146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1803_ u_cpu.cpu.mem_bytecnt\[1\] _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1734_ _1174_ _1183_ _1184_ u_arbiter.o_wb_cpu_adr\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1665_ u_arbiter.i_wb_cpu_dbus_adr\[11\] _1130_ _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3136__CLK net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1596_ _1072_ u_cpu.cpu.state.ibus_cyc _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2468__C _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout74_I net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2217_ _0390_ _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3197_ _0025_ net45 u_cpu.rf_ram.regzero vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2148_ _0266_ _0312_ _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_22_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2079_ _1244_ _0287_ _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2285__I0 u_arbiter.i_wb_cpu_rdt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2512__I1 u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1779__A2 u_cpu.cpu.immdec.imm31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2976__A1 _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_scanchain_local.scan_flop\[52\] u_scanchain_local.module_data_in\[51\] net141 u_arbiter.o_wb_cpu_adr\[14\]
+ net28 u_scanchain_local.module_data_in\[52\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__3159__CLK net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2751__I1 u_arbiter.i_wb_cpu_dbus_adr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3120_ _0144_ net77 u_cpu.cpu.bufreg.lsb\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2900__A1 u_cpu.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3051_ _0076_ net103 u_arbiter.i_wb_cpu_dbus_dat\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2002_ u_cpu.cpu.bufreg.c_r _0227_ _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_64_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2967__A1 _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2904_ _0247_ _0966_ _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_17_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2835_ _0912_ _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2195__A2 _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2766_ u_cpu.cpu.state.o_cnt_r\[1\] _1281_ _1247_ _0257_ _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1717_ _1169_ _1170_ _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2697_ _1288_ _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1648_ u_arbiter.i_wb_cpu_dbus_adr\[8\] _1116_ _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1579_ _1057_ _1054_ _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2661__C _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2186__A2 _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2249__I0 u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2413__A3 _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2620_ _0761_ _0756_ _0762_ _0567_ _0103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_fanout124_I net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2177__A2 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2551_ _0694_ _0700_ _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2482_ u_cpu.cpu.immdec.imm24_20\[1\] _0638_ _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3103_ _0128_ net114 u_arbiter.i_wb_cpu_dbus_adr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3034_ _0059_ net89 u_arbiter.i_wb_cpu_dbus_dat\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout37_I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2762__B _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1612__A1 _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2818_ _1147_ _0899_ _0901_ u_cpu.cpu.ctrl.o_ibus_adr\[17\] _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2749_ u_arbiter.i_wb_cpu_dbus_adr\[25\] u_arbiter.i_wb_cpu_dbus_adr\[26\] _0855_
+ _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2412__I0 u_arbiter.i_wb_cpu_rdt\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2340__A2 _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2991__CLK net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[15\] u_arbiter.i_wb_cpu_rdt\[12\] net130 u_arbiter.i_wb_cpu_dbus_dat\[9\]
+ net16 u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__2867__B1 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.input_buf_clk net1 u_scanchain_local.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_19_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1842__A1 _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1982_ u_cpu.cpu.immdec.imm11_7\[3\] _1387_ _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2642__I0 u_arbiter.i_wb_cpu_rdt\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2603_ _0622_ _0510_ _0748_ _0497_ _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2534_ u_cpu.cpu.immdec.imm30_25\[1\] _0542_ _0685_ _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2465_ _0552_ _0502_ _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2396_ _0542_ _0559_ _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2322__A2 _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2086__A1 _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3017_ _0042_ net70 u_cpu.cpu.ctrl.i_jump vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_3_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2712__S _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2511__I _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[62\]_CLK net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout130 net132 net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout141 net143 net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_93_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2077__A1 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[15\]_CLK net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2421__I _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2001__A1 _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2552__A2 _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2250_ _0414_ _0415_ _0417_ _0418_ _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2577__B _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2181_ _0369_ _0057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2068__A1 _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1965_ _1202_ _1375_ _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2240__A1 _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1896_ _1334_ _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2517_ _0641_ _0669_ _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2448_ _0575_ _0594_ _0455_ _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2379_ _0460_ _0463_ _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_5_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2707__S _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2059__A1 u_cpu.raddr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_cpu.rf_ram.RAM0_WEN[3] net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1806__A1 _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3042__CLK net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3192__CLK net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2534__A2 _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2397__B _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[8\] u_arbiter.i_wb_cpu_rdt\[5\] net137 u_arbiter.i_wb_cpu_dbus_dat\[2\]
+ net24 u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_48_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2470__A1 _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1750_ u_arbiter.i_wb_cpu_dbus_adr\[30\] _1116_ _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1681_ _1140_ _1137_ u_cpu.cpu.ctrl.o_ibus_adr\[15\] _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2151__I _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2302_ _0470_ _0432_ _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2233_ u_arbiter.i_wb_cpu_rdt\[29\] _0318_ _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2164_ _0357_ _0052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_22_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2095_ u_cpu.cpu.bne_or_bge _1028_ _1035_ _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3065__CLK net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2997_ _0010_ net51 u_cpu.rf_ram_if.rdata1\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1948_ _1366_ _0012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1879_ _1048_ _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_66_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2516__A2 _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2664__C _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2452__A1 _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2507__A2 _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2920_ _0975_ _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_u_scanchain_local.scan_flop\[8\]_CLK net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2851_ _0921_ _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2782_ u_arbiter.i_wb_cpu_ibus_adr\[1\] _0877_ _0880_ _1084_ _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1802_ u_cpu.cpu.decode.op22 _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1733_ u_arbiter.i_wb_cpu_dbus_adr\[26\] _1172_ _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1664_ _1089_ _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1595_ net2 _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2216_ _0392_ _0393_ _0068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_fanout67_I net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3196_ _0024_ net45 u_cpu.rf_ram.rdata\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2147_ _0317_ _0343_ _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2682__A1 _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2078_ _0286_ _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2434__A1 _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2285__I1 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2673__A1 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2425__A1 _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[30\]_D u_arbiter.i_wb_cpu_rdt\[27\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_scanchain_local.scan_flop\[45\] u_scanchain_local.module_data_in\[44\] net147 u_arbiter.o_wb_cpu_adr\[7\]
+ net31 u_scanchain_local.module_data_in\[45\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_5_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[16\]_SE net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2900__A2 _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3050_ _0075_ net103 u_arbiter.i_wb_cpu_dbus_dat\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2001_ _1207_ _0223_ _0225_ _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_64_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2664__A1 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2416__A1 _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2903_ _1083_ _0965_ _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_32_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2967__A2 _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2834_ _1169_ _0906_ _0908_ u_cpu.cpu.ctrl.o_ibus_adr\[24\] _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_u_scanchain_local.scan_flop\[23\]_SI u_arbiter.i_wb_cpu_dbus_dat\[17\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3103__CLK net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[21\]_D u_arbiter.i_wb_cpu_rdt\[18\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_2765_ _0864_ _0866_ _0868_ _0233_ _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1716_ u_cpu.cpu.ctrl.o_ibus_adr\[22\] u_cpu.cpu.ctrl.o_ibus_adr\[21\] u_cpu.cpu.ctrl.o_ibus_adr\[20\]
+ _1157_ _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_2696_ _0829_ _0112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1647_ _1089_ _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1578_ _1024_ _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_67_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3179_ _0200_ net67 u_cpu.cpu.genblk3.csr.mcause3_0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2655__A1 u_cpu.cpu.immdec.imm19_12_20\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2407__A1 _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1630__A2 _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[12\]_D u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[39\]_SE net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2894__A1 _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2646__A1 _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2249__I1 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout117_I net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2550_ _0598_ _0697_ _0698_ _0699_ _0537_ _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_12_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2481_ _0411_ _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2885__A1 _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3102_ _0127_ net98 u_arbiter.i_wb_cpu_dbus_adr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3033_ _0058_ net89 u_arbiter.i_wb_cpu_dbus_dat\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2637__A1 _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2817_ _0902_ _0160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2748_ _0858_ _0135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2412__I1 u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2679_ _0590_ u_arbiter.i_wb_cpu_rdt\[19\] _0496_ _0815_ _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_28_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3149__CLK net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2244__I _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2867__A1 _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2867__B2 _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2095__A2 _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1981_ _1385_ _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2642__I1 u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2602_ _0746_ _0747_ _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2533_ _0530_ _0684_ _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2464_ _0621_ _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2395_ _0517_ _0551_ _0558_ _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2858__B2 _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3016_ _0041_ net66 u_cpu.cpu.mem_if.signbit vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_58_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2064__I _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2794__B1 _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout120 net121 net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout131 net132 net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout142 net143 net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_41_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2077__A2 _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1588__A1 _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2180_ u_arbiter.i_wb_cpu_rdt\[12\] _0368_ _0323_ u_arbiter.i_wb_cpu_dbus_dat\[12\]
+ _0361_ u_arbiter.i_wb_cpu_dbus_dat\[13\] _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_120_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2149__I _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1988__I _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1579__A1 _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1964_ _1020_ u_cpu.rf_ram_if.rcnt\[1\] u_cpu.rf_ram_if.rcnt\[2\] _1375_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_105_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2240__A2 u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2612__I _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1895_ u_cpu.rf_ram.rdata\[1\] u_cpu.rf_ram.data\[1\] _1333_ _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout97_I net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2516_ u_cpu.cpu.immdec.imm30_25\[0\] _0476_ _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2447_ _0455_ _0575_ _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2487__C _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2378_ _0513_ _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1806__A2 _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2008__B _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2432__I _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1680_ _1139_ _1142_ u_arbiter.o_wb_cpu_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2588__B _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2301_ _0453_ _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2232_ u_arbiter.i_wb_cpu_dbus_dat\[30\] _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2289__A2 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2163_ u_arbiter.i_wb_cpu_rdt\[7\] _0321_ _0323_ u_arbiter.i_wb_cpu_dbus_dat\[7\]
+ _0352_ u_arbiter.i_wb_cpu_dbus_dat\[8\] _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2094_ _1258_ _1237_ _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_59_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_u_scanchain_local.scan_flop\[61\]_CLK net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout12_I u_arbiter.i_wb_cpu_ack vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2996_ _0009_ net53 u_cpu.rf_ram_if.rdata1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1947_ u_cpu.rf_ram_if.rdata1\[6\] _1365_ u_cpu.rf_ram_if.rtrig1 _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1972__A1 _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1878_ _1314_ _1316_ _1319_ _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2718__S _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[14\]_CLK net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2452__A2 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2252__I _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2427__I _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout147_I net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2850_ u_cpu.cpu.ctrl.o_ibus_adr\[30\] _0876_ _0879_ u_cpu.cpu.ctrl.o_ibus_adr\[31\]
+ _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_54_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2590__C _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1801_ u_cpu.cpu.state.o_cnt_r\[3\] _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_106_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2781_ _0881_ _0145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1732_ _1181_ _1182_ _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_15_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1663_ _1119_ _1112_ _1113_ _1128_ _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1706__A1 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1594_ u_arbiter.i_wb_cpu_ibus_adr\[0\] _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2215_ u_arbiter.i_wb_cpu_rdt\[23\] _0321_ _0351_ u_arbiter.i_wb_cpu_dbus_dat\[23\]
+ _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3032__CLK net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3195_ _0023_ net45 u_cpu.rf_ram.rdata\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2146_ u_arbiter.i_wb_cpu_dbus_dat\[4\] _0259_ _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2682__A2 u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2077_ net2 _1217_ _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2434__A2 _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3182__CLK net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2273__S _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2979_ _1353_ _0024_ _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2800__I _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2956__B _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2673__A2 _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2425__A2 _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[38\] u_scanchain_local.module_data_in\[37\] net137 u_arbiter.o_wb_cpu_adr\[0\]
+ net24 u_scanchain_local.module_data_in\[38\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_5_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3055__CLK net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2361__A1 _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2000_ _1207_ u_cpu.cpu.bufreg.c_r _0223_ _0225_ _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2664__A2 _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2902_ u_arbiter.i_wb_cpu_ack u_arbiter.o_wb_cpu_adr\[1\] _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2833_ _0911_ _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2764_ _0228_ _0231_ _0867_ _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1715_ u_cpu.cpu.ctrl.o_ibus_adr\[23\] _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2695_ u_cpu.cpu.alu.cmp_r _0304_ _1232_ _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1646_ _1112_ _1113_ _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_63_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1577_ u_cpu.cpu.immdec.imm19_12_20\[7\] _1027_ _1055_ u_cpu.cpu.immdec.imm24_20\[3\]
+ _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_63_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2352__A1 _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1950__I1 _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2104__A1 _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3178_ _0199_ net76 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2129_ _0325_ _0327_ _0267_ _0328_ _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2407__A2 _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2591__A1 _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3078__CLK net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[7\]_CLK net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2343__A1 _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1941__I1 _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2906__S _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2480_ _0615_ _0637_ _0088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2334__A1 _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3101_ _0126_ net98 u_arbiter.i_wb_cpu_dbus_adr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1932__I1 _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2885__A2 _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3032_ _0057_ net89 u_arbiter.i_wb_cpu_dbus_dat\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2637__A2 _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2816_ u_cpu.cpu.ctrl.o_ibus_adr\[15\] _0899_ _0901_ _1147_ _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2747_ u_arbiter.i_wb_cpu_dbus_adr\[24\] u_arbiter.i_wb_cpu_dbus_adr\[25\] _0855_
+ _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2678_ _1082_ _0337_ _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2573__A1 _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1629_ u_cpu.cpu.genblk1.align.ctrl_misal u_cpu.cpu.ctrl.o_ibus_adr\[4\] u_cpu.cpu.ctrl.o_ibus_adr\[3\]
+ u_cpu.cpu.ctrl.o_ibus_adr\[2\] _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_67_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2325__A1 _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2628__A2 _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[0\]_SE net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2564__A1 _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2260__I _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2867__A2 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1604__I _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2619__A2 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1980_ _1065_ _1380_ _1385_ _1386_ u_cpu.rf_ram.addr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2601_ _0579_ _0442_ _0548_ _0621_ _0583_ _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__2555__A1 _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2532_ _1232_ _0683_ _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2463_ _0418_ _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2394_ _0553_ _0555_ _0557_ _0434_ _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1905__I1 u_cpu.rf_ram.data\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2546__S _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3015_ _0040_ net70 u_cpu.cpu.state.genblk1.misalign_trap_sync_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout42_I net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout121 net122 net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout110 net123 net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout143 net149 net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout132 net133 net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_41_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2234__B1 _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1588__A2 _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2001__A3 _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xu_scanchain_local.scan_flop\[20\] u_arbiter.i_wb_cpu_rdt\[17\] net127 u_arbiter.i_wb_cpu_dbus_dat\[14\]
+ net13 u_arbiter.i_wb_cpu_rdt\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2170__C1 _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2165__I _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1963_ _1374_ _0006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1894_ _1203_ _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_18_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3139__CLK net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2515_ _0498_ _0663_ _0667_ _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2446_ _0251_ u_arbiter.i_wb_cpu_rdt\[4\] _0604_ _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_142_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2377_ _1235_ _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1806__A3 _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2803__I _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1990__A2 _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2914__S _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[68\] u_scanchain_local.module_data_in\[67\] net147 u_arbiter.o_wb_cpu_adr\[30\]
+ net32 u_scanchain_local.module_data_in\[68\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_102_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2869__B _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1733__A2 _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2300_ _0465_ _0468_ _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2231_ u_arbiter.i_wb_cpu_dbus_dat\[29\] _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2162_ _0355_ _0356_ _0051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2093_ _1321_ _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_4_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2995_ _0008_ net53 u_cpu.rf_ram_if.rdata1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1946_ _1352_ _0023_ _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_30_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1877_ _1316_ _1318_ _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1972__A2 _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1724__A2 _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2429_ _1081_ _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__1903__S _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2988__A1 _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2734__S _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1800_ _1215_ _1216_ _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2780_ _1071_ _0877_ _0880_ u_arbiter.i_wb_cpu_ibus_adr\[1\] _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_12_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1731_ u_cpu.cpu.ctrl.o_ibus_adr\[25\] u_cpu.cpu.ctrl.o_ibus_adr\[24\] u_cpu.cpu.ctrl.o_ibus_adr\[23\]
+ _1170_ _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_8_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1662_ u_cpu.cpu.ctrl.o_ibus_adr\[11\] u_cpu.cpu.ctrl.o_ibus_adr\[10\] _1128_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2903__A1 _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1593_ _1027_ u_cpu.rf_ram_if.wtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2214_ u_arbiter.i_wb_cpu_dbus_dat\[24\] _0352_ _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3194_ _0022_ net46 u_cpu.rf_ram.rdata\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2145_ _0337_ _0339_ _0341_ _0342_ _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2076_ _0247_ _0285_ _0035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1678__B _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2978_ _0877_ _1012_ _1013_ _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1929_ _1352_ _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2370__A2 _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2830__B1 _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[60\]_CLK net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2361__A2 _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1624__A1 _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2901_ _0728_ _0964_ _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2416__A3 _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[62\]_SE net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2173__I _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2832_ u_cpu.cpu.ctrl.o_ibus_adr\[22\] _0906_ _0908_ _1169_ _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2763_ _0228_ _0231_ _0243_ _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1714_ _1132_ _1167_ _1168_ u_arbiter.o_wb_cpu_adr\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_u_scanchain_local.scan_flop\[13\]_CLK net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2694_ _0826_ _0827_ _0828_ _0111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1645_ _1112_ _1113_ _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[28\]_CLK net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1576_ _1023_ _1054_ _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA_fanout72_I net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2348__I _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3177_ _0198_ net92 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2128_ net39 _0316_ _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2059_ u_cpu.raddr\[0\] _0272_ _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_74_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2591__A2 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2718__I1 u_arbiter.i_wb_cpu_dbus_adr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2343__A2 _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2894__A3 _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[50\] u_scanchain_local.module_data_in\[49\] net141 u_arbiter.o_wb_cpu_adr\[12\]
+ net27 u_scanchain_local.module_data_in\[50\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_51_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2582__A2 _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3172__CLK net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2334__A2 _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3100_ _0125_ net98 u_arbiter.i_wb_cpu_dbus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3031_ _0056_ net93 u_arbiter.i_wb_cpu_dbus_dat\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2270__A1 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2815_ _0879_ _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2746_ _0857_ _0134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2677_ _0562_ _0619_ _0576_ _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1628_ u_cpu.cpu.ctrl.o_ibus_adr\[5\] _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1559_ _1029_ u_cpu.cpu.decode.op21 _1034_ _1037_ _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__1911__S _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2089__A1 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2027__B _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3045__CLK net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3195__CLK net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2013__A1 _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2564__A2 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2917__S _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1827__A1 u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1620__I _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout122_I net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2600_ _0470_ _0738_ _0745_ _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2531_ _0297_ _0682_ _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2462_ _0553_ _0619_ _0456_ _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_87_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2400__B _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2393_ _0556_ _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1818__A1 _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3014_ _0039_ net79 u_cpu.cpu.state.o_cnt_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3068__CLK net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2491__A1 _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout35_I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[6\]_CLK net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2794__A2 _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2729_ u_arbiter.i_wb_cpu_dbus_adr\[16\] u_arbiter.i_wb_cpu_dbus_adr\[17\] _0843_
+ _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout111 net113 net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout122 net123 net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout100 net124 net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_114_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout144 net149 net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout133 net134 net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_80_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1809__A1 _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2537__A2 _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1615__I _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[13\] u_arbiter.i_wb_cpu_rdt\[10\] net130 u_arbiter.i_wb_cpu_dbus_dat\[7\]
+ net16 u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_2_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1899__I1 u_cpu.rf_ram.data\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2170__B1 _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3210__CLK net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2890__B _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2225__A1 u_arbiter.i_wb_cpu_rdt\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1962_ u_cpu.rf_ram_if.rdata0\[7\] _1365_ _1057_ _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1893_ _1210_ _1213_ _0017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2514_ _0592_ _0539_ _0598_ _0666_ _0508_ _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_2445_ _1080_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[4\] _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_64_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2161__B1 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2376_ _0450_ _0538_ _0511_ _0539_ _0540_ _0081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_72_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_cpu.rf_ram.RAM0_WEN[0] net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1806__A4 _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2767__A2 _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1990__A3 _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2152__B1 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2455__A1 _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2455__B2 _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2930__S _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[19\]_SE net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2230_ _0402_ _0073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2161_ u_arbiter.i_wb_cpu_rdt\[6\] _0339_ _0348_ u_arbiter.i_wb_cpu_dbus_dat\[6\]
+ _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_47_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2092_ u_cpu.cpu.ctrl.i_jump _0287_ _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2446__A1 _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2994_ _0007_ net53 u_cpu.rf_ram_if.rdata1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3106__CLK net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1945_ _1364_ _0011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1876_ _1317_ u_arbiter.i_wb_cpu_dbus_dat\[8\] u_arbiter.i_wb_cpu_dbus_dat\[16\]
+ u_arbiter.i_wb_cpu_dbus_dat\[24\] u_cpu.cpu.bufreg.lsb\[0\] _1026_ _1318_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_31_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2428_ _0510_ _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2359_ _0521_ _0524_ _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2437__A1 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2035__B _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[6\] u_arbiter.i_wb_cpu_rdt\[3\] net136 u_arbiter.i_wb_cpu_dbus_dat\[0\]
+ net21 u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_76_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2925__S _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3129__CLK net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[33\]_D u_arbiter.i_wb_cpu_rdt\[30\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1730_ u_cpu.cpu.ctrl.o_ibus_adr\[26\] _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2600__A1 _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1661_ _1124_ _1120_ u_cpu.cpu.ctrl.o_ibus_adr\[11\] _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2599__C _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1592_ _1060_ _1070_ _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2213_ _0391_ _0067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_61_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1803__I u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3193_ _0021_ net44 u_cpu.rf_ram.rdata\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2144_ u_arbiter.i_wb_cpu_dbus_dat\[3\] _0333_ _0338_ _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_82_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2419__A1 _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2075_ _1246_ _0284_ _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_50_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[24\]_D u_arbiter.i_wb_cpu_rdt\[21\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2977_ u_cpu.cpu.state.ibus_cyc _1012_ _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_10_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1928_ u_cpu.rf_ram.regzero _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1859_ _1042_ _1300_ _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1633__A2 _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_u_scanchain_local.scan_flop\[15\]_D u_arbiter.i_wb_cpu_rdt\[12\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2897__A1 _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2361__A3 _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2649__A1 _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2900_ u_cpu.cpu.bufreg.i_sh_signed _0413_ _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2831_ _0910_ _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2762_ u_cpu.cpu.bufreg.i_sh_signed _0243_ _0233_ _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1713_ u_arbiter.i_wb_cpu_dbus_adr\[22\] _1109_ _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2403__B _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2693_ u_cpu.cpu.genblk3.csr.mie_mtie u_cpu.cpu.genblk3.csr.mstatus_mie u_cpu.cpu.genblk3.csr.i_mtip
+ _0827_ _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_67_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1644_ u_cpu.cpu.ctrl.o_ibus_adr\[7\] u_cpu.cpu.ctrl.o_ibus_adr\[6\] u_cpu.cpu.ctrl.o_ibus_adr\[5\]
+ _1101_ _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__2888__A1 u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1575_ _1038_ _1053_ _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3176_ _0197_ net76 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout65_I net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2127_ _0313_ _0326_ _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1863__A2 _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2058_ u_cpu.raddr\[0\] _0272_ _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2040__A2 _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2591__A3 _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1926__I0 u_cpu.rf_ram_if.wdata1_r\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[43\] u_scanchain_local.module_data_in\[42\] net138 u_arbiter.o_wb_cpu_adr\[5\]
+ net23 u_scanchain_local.module_data_in\[43\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3030_ _0055_ net93 u_arbiter.i_wb_cpu_dbus_dat\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2814_ _0900_ _0159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_121_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2745_ u_arbiter.i_wb_cpu_dbus_adr\[23\] u_arbiter.i_wb_cpu_dbus_adr\[24\] _0855_
+ _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_133_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2676_ _0781_ _0811_ _0812_ _0813_ _0108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_114_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1627_ _1094_ _1098_ _1099_ u_arbiter.o_wb_cpu_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1972__B _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1781__A1 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1558_ _1036_ _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_115_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2089__A2 _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3159_ _0180_ net60 u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2013__A2 _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2564__A3 _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[52\]_SE net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[12\]_CLK net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_u_scanchain_local.scan_flop\[27\]_CLK net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout115_I net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2530_ _1320_ _1265_ _1204_ _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2461_ _0618_ _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2392_ _0479_ _0457_ _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_25_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3215__D u_cpu.rf_ram_if.wdata1_r\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3013_ _0038_ net80 u_cpu.cpu.state.o_cnt_r\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1818__A2 _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout28_I net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2728_ _0847_ _0126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1754__A1 _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2659_ _0576_ _0618_ _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfanout112 net113 net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout101 net104 net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
Xfanout145 net146 net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout134 net151 net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout123 net124 net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_86_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3012__CLK net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1721__I _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2482__A2 _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2753__S _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2234__A2 _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1993__A1 u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2501__B _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2928__S _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2170__A1 u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2225__A2 _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1961_ _1373_ _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1892_ _1298_ _1332_ u_cpu.cpu.o_wdata0 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2513_ _0414_ _0528_ _0664_ _0665_ _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2411__B _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2444_ _0471_ _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3035__CLK net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2375_ _1266_ _0514_ _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2161__A1 u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2161__B2 u_arbiter.i_wb_cpu_dbus_dat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3185__CLK net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1975__A1 u_cpu.cpu.decode.op26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1917__S _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2152__A1 u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2455__A2 _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1966__A1 u_cpu.raddr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3058__CLK net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2391__A1 _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2160_ u_arbiter.i_wb_cpu_dbus_dat\[7\] _0354_ _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2091_ _0294_ _0295_ _0040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2446__A2 u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2993_ _0031_ net64 u_cpu.raddr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1944_ u_cpu.rf_ram_if.rdata1\[5\] _1363_ _1355_ _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1875_ u_arbiter.i_wb_cpu_dbus_dat\[0\] _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout95_I net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2427_ _0514_ _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2134__A1 _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2358_ _0523_ _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2685__A2 _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2289_ _0446_ _0457_ _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_42_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3200__CLK net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2051__B _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2373__A1 _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2125__A1 u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1660_ _1123_ _1126_ u_arbiter.o_wb_cpu_adr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1591_ _1064_ _1065_ _1069_ _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2212_ u_arbiter.i_wb_cpu_rdt\[22\] _0368_ _0390_ u_arbiter.i_wb_cpu_dbus_dat\[22\]
+ _0361_ u_arbiter.i_wb_cpu_dbus_dat\[23\] _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_61_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3192_ _0020_ net46 u_cpu.rf_ram.rdata\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2143_ u_arbiter.i_wb_cpu_dbus_dat\[4\] _0317_ _0313_ _0340_ _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1890__A3 _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2074_ _1315_ _0281_ _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2136__B _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2976_ _0412_ _0286_ _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout10_I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1927_ _1351_ u_cpu.rf_ram.i_wdata\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1858_ _1299_ _1206_ _1226_ _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__2355__A1 _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1789_ _1206_ _1229_ _1232_ _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_44_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2107__A1 _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[3\]_SE net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2046__B _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2830__A2 _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2594__A1 _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2897__A2 _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2936__S _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2830_ u_cpu.cpu.ctrl.o_ibus_adr\[21\] _0906_ _0908_ u_cpu.cpu.ctrl.o_ibus_adr\[22\]
+ _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_fanout145_I net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2761_ _0864_ _0233_ _0865_ _0141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1712_ u_cpu.cpu.ctrl.o_ibus_adr\[22\] _1166_ _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2585__A1 u_cpu.cpu.immdec.imm31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2692_ _0277_ _0243_ _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1643_ u_cpu.cpu.ctrl.o_ibus_adr\[8\] _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__2403__C _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3218__D u_cpu.rf_ram_if.wdata1_r\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2337__A1 _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2888__A2 _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1574_ _1044_ _1052_ _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1935__I1 _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3175_ _0196_ net92 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2126_ _1317_ net39 _0314_ _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout58_I net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2057_ _1375_ _0270_ _0272_ _0029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_63_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2959_ _0277_ _1262_ _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2380__I _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2328__A1 _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2879__A2 _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3119__CLK net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1926__I1 u_cpu.cpu.o_wdata0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2500__A1 _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2567__A1 _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xu_scanchain_local.scan_flop\[36\] u_scanchain_local.module_data_in\[35\] net144 u_arbiter.i_wb_cpu_dbus_dat\[30\]
+ net30 u_scanchain_local.module_data_in\[36\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__1917__I1 u_cpu.rf_ram_if.wdata1_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2813_ _1140_ _0899_ _0894_ u_cpu.cpu.ctrl.o_ibus_adr\[15\] _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2744_ _0856_ _0133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2675_ u_cpu.cpu.immdec.imm19_12_20\[7\] _0755_ _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1626_ u_arbiter.i_wb_cpu_dbus_adr\[4\] _1091_ _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1781__A2 _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1557_ _1035_ u_cpu.cpu.bne_or_bge _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2576__S _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3158_ _0179_ net60 u_cpu.cpu.immdec.imm11_7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2109_ u_cpu.cpu.bufreg.lsb\[1\] u_cpu.cpu.mem_bytecnt\[1\] _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3089_ _0114_ net106 u_arbiter.i_wb_cpu_dbus_adr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2549__A1 _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1772__A2 _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3091__CLK net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1827__A3 _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2237__B1 _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout108_I net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2460_ _0617_ _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2391_ _0554_ _0468_ _0509_ _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3012_ _0037_ net79 u_cpu.cpu.state.o_cnt_r\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2144__B _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2727_ u_arbiter.i_wb_cpu_dbus_adr\[15\] u_arbiter.i_wb_cpu_dbus_adr\[16\] _0843_
+ _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2251__I0 u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2951__A1 _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2658_ u_arbiter.i_wb_cpu_rdt\[17\] u_arbiter.i_wb_cpu_rdt\[1\] _1081_ _0797_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xfanout113 net116 net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout102 net104 net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1609_ u_cpu.cpu.ctrl.o_ibus_adr\[2\] _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2589_ _0728_ _0729_ _0735_ _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_102_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout146 net148 net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout124 net125 net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout135 net140 net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_68_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2219__B1 _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1993__A2 _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1745__A2 _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2942__B2 _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2501__C _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2170__A2 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1912__I _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1960_ u_cpu.rf_ram_if.rdata0\[6\] _1363_ _1057_ _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_15_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1891_ _1066_ _1331_ _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2512_ u_arbiter.i_wb_cpu_rdt\[24\] u_arbiter.i_wb_cpu_rdt\[8\] _1082_ _0665_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2443_ u_arbiter.i_wb_cpu_rdt\[22\] u_arbiter.i_wb_cpu_rdt\[6\] _1081_ _0602_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2374_ _0436_ _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2161__A2 _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1822__I _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_75_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[42\]_SE net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1975__A2 u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[11\]_CLK net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[26\]_CLK net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2152__A2 _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2997__CLK net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1642__I _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2090_ _0217_ _0220_ _0032_ _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_111_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[65\]_SE net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1654__A1 _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2992_ _0030_ net63 u_cpu.raddr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1943_ _1352_ _0022_ _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_119_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1874_ _1236_ _1246_ _1315_ _1037_ _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1709__A2 _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3002__CLK net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2757__I1 u_arbiter.i_wb_cpu_dbus_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1590__B1 _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2426_ _1039_ _0515_ _0586_ _0085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3152__CLK net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout88_I net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2357_ _0250_ u_arbiter.i_wb_cpu_rdt\[10\] _0522_ _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2288_ _0447_ _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2070__A1 _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2332__B _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2051__C _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xu_scanchain_local.scan_flop\[66\] u_scanchain_local.module_data_in\[65\] net145 u_arbiter.o_wb_cpu_adr\[28\]
+ net33 u_scanchain_local.module_data_in\[66\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__3025__CLK net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1590_ u_cpu.cpu.csr_imm _1023_ _1055_ u_cpu.cpu.immdec.imm24_20\[0\] _1068_ _1069_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_67_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2211_ _0322_ _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3191_ _0019_ net46 u_cpu.rf_ram.rdata\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2142_ _0317_ _0259_ _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2073_ _1315_ _0281_ _0283_ _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1627__A1 _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2052__A1 u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2975_ _0246_ u_cpu.cpu.genblk3.csr.timer_irq_r _0828_ _1011_ _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_33_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1926_ u_cpu.rf_ram_if.wdata1_r\[7\] u_cpu.cpu.o_wdata0 _1350_ _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1857_ u_cpu.cpu.alu.i_rs1 u_cpu.cpu.alu.add_cy_r _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2355__A2 u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1788_ _1231_ _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_131_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2409_ _0466_ _0472_ _0570_ _0517_ _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_130_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2378__I _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3048__CLK net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2594__A2 u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2806__B1 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2282__A1 _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_fanout138_I net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2034__A1 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2760_ u_arbiter.i_wb_cpu_dbus_adr\[30\] _0233_ _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1711_ u_cpu.cpu.ctrl.o_ibus_adr\[21\] _1160_ _1157_ _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2691_ u_cpu.cpu.genblk3.csr.timer_irq_r _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1642_ _1090_ _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2337__A2 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1573_ _1046_ _1051_ _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3174_ _0195_ net91 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2125_ u_arbiter.i_wb_cpu_dbus_dat\[2\] _0314_ _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2056_ _0271_ _1021_ _1022_ _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_41_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2025__A1 _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2958_ _0997_ _0998_ _0999_ _1261_ _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1909_ u_cpu.rf_ram_if.genblk1.wtrig0_r _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_68_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2889_ _0592_ _0484_ _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2328__A2 _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1941__S _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2836__I _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2504__C _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2567__A2 u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[29\] u_arbiter.i_wb_cpu_rdt\[26\] net131 u_arbiter.i_wb_cpu_dbus_dat\[23\]
+ net17 u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XANTENNA__3054__D _0079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3213__CLK net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2812_ _0875_ _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2743_ u_arbiter.i_wb_cpu_dbus_adr\[22\] u_arbiter.i_wb_cpu_dbus_adr\[23\] _0855_
+ _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2674_ u_cpu.cpu.immdec.imm19_12_20\[8\] _0568_ _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1625_ u_cpu.cpu.ctrl.o_ibus_adr\[4\] _1097_ _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_126_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1556_ u_cpu.cpu.decode.co_mem_word _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2191__B1 _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_fanout70_I net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1560__I u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2494__B2 _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3157_ _0178_ net61 u_cpu.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2108_ u_cpu.cpu.bufreg.lsb\[1\] u_cpu.cpu.mem_bytecnt\[1\] u_cpu.cpu.mem_bytecnt\[0\]
+ u_cpu.cpu.bufreg.lsb\[0\] _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3088_ _0113_ net105 u_arbiter.i_wb_cpu_dbus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2039_ _1236_ _1048_ _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2549__A2 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2390_ _0516_ _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3011_ _0036_ net79 u_cpu.cpu.state.o_cnt_r\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2476__A1 _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3109__CLK net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2726_ _0846_ _0125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2251__I1 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2400__A1 _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2951__A2 _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2657_ _0781_ _0794_ _0795_ _0796_ _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1608_ _1082_ _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout103 net104 net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_2588_ u_cpu.cpu.immdec.imm7 _0225_ _0690_ _0734_ _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_114_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout114 net116 net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout147 net149 net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout125 net126 net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout136 net140 net136 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1539_ u_cpu.rf_ram_if.rcnt\[0\] _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_41_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3209_ _0213_ net68 u_cpu.rf_ram_if.rgnt vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1690__A2 _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2219__A1 u_arbiter.i_wb_cpu_rdt\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2942__A2 _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[3\]_D u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1890_ _1257_ _1312_ _1313_ _1330_ _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_18_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout120_I net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2394__B1 _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2511_ _0506_ _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2442_ _1040_ _0587_ _0601_ _0086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_64_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2373_ _0533_ _0535_ _0537_ _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_68_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1672__A2 _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout33_I net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1994__B _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1975__A3 _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2709_ _0830_ _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2688__A1 _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2860__A1 _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2376__B1 _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2679__A1 _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xu_scanchain_local.scan_flop\[11\] u_arbiter.i_wb_cpu_rdt\[8\] net134 u_arbiter.i_wb_cpu_dbus_dat\[5\]
+ net20 u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_4_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2991_ _0029_ net63 u_cpu.rf_ram_if.rcnt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1942_ _1362_ _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2603__A1 _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1873_ u_cpu.cpu.mem_bytecnt\[0\] _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_70_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2425_ _0510_ _0573_ _0577_ _0585_ _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__1590__B2 u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1590__A1 u_cpu.cpu.csr_imm vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2356_ _0427_ u_cpu.cpu.genblk1.align.ibus_rdt_concat\[10\] _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_85_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2287_ _0455_ _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_42_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1645__A2 _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[27\]_D u_arbiter.i_wb_cpu_rdt\[24\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2613__B _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1944__S _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2839__I _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xu_cpu.rf_ram.RAM0_152 net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2381__I0 u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1884__A2 u_cpu.cpu.ctrl.i_iscomp vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1636__A2 _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[18\]_D u_arbiter.i_wb_cpu_rdt\[15\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xu_scanchain_local.scan_flop\[59\] u_scanchain_local.module_data_in\[58\] net146 u_arbiter.o_wb_cpu_adr\[21\]
+ net34 u_scanchain_local.module_data_in\[59\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_8_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1572__A1 _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2210_ _0388_ _0389_ _0066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[32\]_SE net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3190_ _0018_ net46 u_cpu.rf_ram.rdata\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2141_ _0338_ _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2072_ _1315_ _0281_ _0282_ _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_u_scanchain_local.scan_flop\[10\]_CLK net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2974_ _1047_ _0287_ _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_u_scanchain_local.scan_flop\[25\]_CLK net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1925_ u_cpu.rf_ram_if.genblk1.wtrig0_r _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_107_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1856_ _1266_ _1280_ _1297_ _1052_ _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1787_ _1230_ _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1563__A1 _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2408_ _0441_ _0543_ _0519_ _0569_ _0564_ _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_2339_ _0480_ _0493_ _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_40_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1866__A2 _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[55\]_SE net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[4\] u_arbiter.i_wb_cpu_rdt\[1\] net135 u_arbiter.i_wb_cpu_dbus_sel\[2\]
+ net22 u_arbiter.i_wb_cpu_rdt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_21_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2034__A2 _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1710_ _1132_ _1164_ _1165_ u_arbiter.o_wb_cpu_adr\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2690_ _0825_ _0110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_126_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1641_ _1094_ _1108_ _1110_ u_arbiter.o_wb_cpu_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2337__A3 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1572_ _1047_ _1050_ _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input5_I io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3173_ _0194_ net91 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2124_ _0316_ _0319_ _0324_ _0045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1848__A2 u_cpu.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2055_ _1020_ _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_63_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2957_ _1047_ _0998_ _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1908_ _1340_ _0024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2888_ u_cpu.cpu.immdec.imm11_7\[3\] _0930_ _0953_ _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1784__A1 _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1839_ u_cpu.cpu.state.o_cnt_r\[0\] _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2389__I _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3015__CLK net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3165__CLK net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout150_I net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2811_ _0898_ _0158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_34_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2742_ _1288_ _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_30_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1766__A1 u_cpu.rf_ram.data\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2673_ _0529_ _0806_ _0810_ _0412_ _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_126_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1624_ _1083_ u_cpu.cpu.ctrl.o_ibus_adr\[3\] _1084_ _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__3038__CLK net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1555_ _1030_ _1033_ _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_28_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2191__A1 u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout63_I net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2494__A2 _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3188__CLK net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3156_ _0177_ net49 u_cpu.cpu.immdec.imm11_7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3087_ _0112_ net65 u_cpu.cpu.alu.cmp_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2107_ _0247_ _0278_ _0308_ _0044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2038_ _0247_ _0255_ _0027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1952__S u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2237__A2 _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xu_scanchain_local.scan_flop\[41\] u_scanchain_local.module_data_in\[40\] net138 u_arbiter.o_wb_cpu_adr\[3\]
+ net23 u_scanchain_local.module_data_in\[41\] vdd vss gf180mcu_fd_sc_mcu7t5v0__sdffq_1
XFILLER_108_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2476__A2 _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3010_ _0035_ net69 u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2725_ u_arbiter.i_wb_cpu_dbus_adr\[14\] u_arbiter.i_wb_cpu_dbus_adr\[15\] _0843_
+ _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2400__A2 _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2656_ u_cpu.cpu.immdec.imm19_12_20\[5\] _0781_ _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1607_ _1081_ _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout104 net110 net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_2587_ _0730_ _0731_ _0733_ _0225_ _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xfanout115 net116 net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout137 net139 net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout126 net5 net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout148 net149 net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_45_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3208_ _0212_ net50 u_cpu.rf_ram_if.rdata0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3139_ _0161_ net98 u_cpu.cpu.ctrl.o_ibus_adr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2219__A2 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2616__B _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1978__A1 _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3203__CLK net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout113_I net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2394__B2 _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2394__A1 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2510_ _0539_ _0527_ _0651_ _0662_ _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_143_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2441_ _0588_ _0591_ _0597_ _0600_ _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2372_ _0536_ _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2449__A2 _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout26_I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2708_ _0836_ _0117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2385__A1 _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2137__A1 u_arbiter.i_wb_cpu_rdt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2639_ u_cpu.cpu.immdec.imm19_12_20\[5\] _0489_ _0755_ _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2932__I0 u_arbiter.i_wb_cpu_rdt\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_u_scanchain_local.scan_flop\[6\]_SE net136 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1663__A3 _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2376__B2 _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2679__A2 u_arbiter.i_wb_cpu_rdt\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2923__I0 u_arbiter.i_wb_cpu_rdt\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2300__A1 _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2990_ _0028_ net53 u_cpu.rf_ram_if.rcnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1941_ u_cpu.rf_ram_if.rdata1\[4\] _1361_ _1355_ _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2603__A2 _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1872_ u_cpu.cpu.mem_if.signbit _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_30_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2367__A1 _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2119__A1 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2424_ _0530_ _0508_ _0581_ _0584_ _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_142_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1590__A2 _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2914__I0 u_arbiter.i_wb_cpu_rdt\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2355_ _0430_ u_arbiter.i_wb_cpu_rdt\[11\] _0520_ _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2286_ _0453_ _0454_ _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2070__A3 _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1956__I1 _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1581__A2 _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2530__A1 _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1960__S _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3071__CLK net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2521__A1 _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2140_ _0320_ _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2071_ _1072_ _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2973_ _0537_ _1010_ _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1924_ _1349_ u_cpu.rf_ram.i_wdata\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2052__A3 _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1855_ _1265_ _1296_ _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1786_ u_cpu.cpu.state.o_cnt_r\[1\] u_cpu.cpu.state.o_cnt_r\[0\] u_cpu.cpu.state.o_cnt_r\[3\]
+ u_cpu.cpu.state.o_cnt_r\[2\] _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA__1938__I1 _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2760__A1 u_arbiter.i_wb_cpu_dbus_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout93_I net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1563__A2 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2407_ _0539_ _0438_ _0525_ _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_58_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2338_ _0411_ _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2269_ _0430_ u_arbiter.i_wb_cpu_rdt\[5\] _0437_ _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2579__A1 _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3094__CLK net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2200__B1 _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2503__A1 _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2806__A2 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2290__I0 u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1640_ u_arbiter.i_wb_cpu_dbus_adr\[7\] _1109_ _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1571_ u_cpu.cpu.decode.op21 _1049_ _1042_ _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__1664__I _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3172_ _0193_ net91 u_cpu.cpu.genblk1.align.ibus_rdt_concat\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2123_ u_arbiter.i_wb_cpu_rdt\[0\] _0321_ _0323_ _1317_ _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2054_ _1020_ _0270_ _0028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_63_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2956_ _0277_ _1253_ _1262_ _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1907_ u_cpu.rf_ram.rdata\[7\] u_cpu.rf_ram.data\[7\] net8 _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2887_ _1389_ _0930_ _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1838_ _1267_ _1279_ _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2981__A1 _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1769_ _1211_ _1212_ u_cpu.rf_ram.rdata\[0\] _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_106_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2619__B _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_u_scanchain_local.scan_flop\[22\]_SE net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2272__I0 u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2972__A1 u_cpu.cpu.ctrl.i_iscomp vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput6 net6 io_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_141_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_u_scanchain_local.scan_flop\[24\]_CLK net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_u_scanchain_local.scan_flop\[39\]_CLK net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2810_ u_cpu.cpu.ctrl.o_ibus_adr\[13\] _0892_ _0894_ _1140_ _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_fanout143_I net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2741_ _0854_ _0132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2963__A1 u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2672_ _0466_ _0799_ _0809_ _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xu_scanchain_local.output_buffers\[3\] net24 u_scanchain_local.clk_out vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1623_ _1094_ _1095_ _1096_ u_arbiter.o_wb_cpu_adr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1554_ _1032_ _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2191__A2 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
.ends

