// This is the unpowered netlist.
module tiny_user_project (user_clock2,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    user_irq,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input user_clock2;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [63:0] la_data_in;
 output [63:0] la_data_out;
 input [63:0] la_oenb;
 output [2:0] user_irq;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire net9;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net10;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net11;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net47;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net48;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net49;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net83;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net84;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net85;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net86;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net87;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net88;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire \mod.timer_irq ;
 wire \mod.u_arbiter.i_wb_cpu_ack ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[10] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[11] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[12] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[13] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[14] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[15] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[16] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[17] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[18] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[19] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[20] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[21] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[22] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[23] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[24] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[25] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[26] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[27] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[28] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[29] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[2] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[30] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[31] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[3] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[4] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[5] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[6] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[7] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[8] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[9] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[0] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[10] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[11] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[12] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[13] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[14] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[15] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[16] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[17] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[18] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[19] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[1] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[20] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[21] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[22] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[23] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[24] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[25] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[26] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[27] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[28] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[29] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[2] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[30] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[31] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[3] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[4] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[5] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[6] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[7] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[8] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[9] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_we ;
 wire \mod.u_arbiter.i_wb_cpu_ibus_adr[0] ;
 wire \mod.u_arbiter.i_wb_cpu_ibus_adr[1] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[0] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[10] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[11] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[12] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[13] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[14] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[15] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[16] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[17] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[18] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[19] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[1] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[20] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[21] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[22] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[23] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[24] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[25] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[26] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[27] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[28] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[29] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[2] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[30] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[31] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[3] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[4] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[5] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[6] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[7] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[8] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[9] ;
 wire \mod.u_cpu.cpu.alu.add_cy_r ;
 wire \mod.u_cpu.cpu.alu.cmp_r ;
 wire \mod.u_cpu.cpu.alu.i_rs1 ;
 wire \mod.u_cpu.cpu.bne_or_bge ;
 wire \mod.u_cpu.cpu.branch_op ;
 wire \mod.u_cpu.cpu.bufreg.c_r ;
 wire \mod.u_cpu.cpu.bufreg.i_sh_signed ;
 wire \mod.u_cpu.cpu.bufreg.lsb[0] ;
 wire \mod.u_cpu.cpu.bufreg.lsb[1] ;
 wire \mod.u_cpu.cpu.bufreg2.i_cnt_done ;
 wire \mod.u_cpu.cpu.csr_d_sel ;
 wire \mod.u_cpu.cpu.csr_imm ;
 wire \mod.u_cpu.cpu.ctrl.i_iscomp ;
 wire \mod.u_cpu.cpu.ctrl.i_jump ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[10] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[11] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[12] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[13] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[14] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[15] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[16] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[17] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[18] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[19] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[20] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[21] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[22] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[23] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[24] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[25] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[26] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[27] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[28] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[29] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[2] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[30] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[31] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[3] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[4] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[5] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[6] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[7] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[8] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[9] ;
 wire \mod.u_cpu.cpu.ctrl.pc_plus_4_cy_r ;
 wire \mod.u_cpu.cpu.ctrl.pc_plus_offset_cy_r ;
 wire \mod.u_cpu.cpu.decode.co_ebreak ;
 wire \mod.u_cpu.cpu.decode.co_mem_word ;
 wire \mod.u_cpu.cpu.decode.op21 ;
 wire \mod.u_cpu.cpu.decode.op22 ;
 wire \mod.u_cpu.cpu.decode.op26 ;
 wire \mod.u_cpu.cpu.decode.opcode[0] ;
 wire \mod.u_cpu.cpu.decode.opcode[1] ;
 wire \mod.u_cpu.cpu.decode.opcode[2] ;
 wire \mod.u_cpu.cpu.genblk1.align.ctrl_misal ;
 wire \mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ;
 wire \mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[10] ;
 wire \mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[11] ;
 wire \mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ;
 wire \mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ;
 wire \mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ;
 wire \mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ;
 wire \mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ;
 wire \mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[2] ;
 wire \mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[3] ;
 wire \mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ;
 wire \mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ;
 wire \mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ;
 wire \mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ;
 wire \mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ;
 wire \mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ;
 wire \mod.u_cpu.cpu.genblk3.csr.mcause31 ;
 wire \mod.u_cpu.cpu.genblk3.csr.mcause3_0[0] ;
 wire \mod.u_cpu.cpu.genblk3.csr.mcause3_0[1] ;
 wire \mod.u_cpu.cpu.genblk3.csr.mcause3_0[2] ;
 wire \mod.u_cpu.cpu.genblk3.csr.mcause3_0[3] ;
 wire \mod.u_cpu.cpu.genblk3.csr.mie_mtie ;
 wire \mod.u_cpu.cpu.genblk3.csr.mstatus_mie ;
 wire \mod.u_cpu.cpu.genblk3.csr.mstatus_mpie ;
 wire \mod.u_cpu.cpu.genblk3.csr.o_new_irq ;
 wire \mod.u_cpu.cpu.genblk3.csr.timer_irq_r ;
 wire \mod.u_cpu.cpu.immdec.imm11_7[0] ;
 wire \mod.u_cpu.cpu.immdec.imm11_7[1] ;
 wire \mod.u_cpu.cpu.immdec.imm11_7[2] ;
 wire \mod.u_cpu.cpu.immdec.imm11_7[3] ;
 wire \mod.u_cpu.cpu.immdec.imm11_7[4] ;
 wire \mod.u_cpu.cpu.immdec.imm19_12_20[0] ;
 wire \mod.u_cpu.cpu.immdec.imm19_12_20[1] ;
 wire \mod.u_cpu.cpu.immdec.imm19_12_20[2] ;
 wire \mod.u_cpu.cpu.immdec.imm19_12_20[3] ;
 wire \mod.u_cpu.cpu.immdec.imm19_12_20[5] ;
 wire \mod.u_cpu.cpu.immdec.imm19_12_20[6] ;
 wire \mod.u_cpu.cpu.immdec.imm19_12_20[7] ;
 wire \mod.u_cpu.cpu.immdec.imm19_12_20[8] ;
 wire \mod.u_cpu.cpu.immdec.imm24_20[0] ;
 wire \mod.u_cpu.cpu.immdec.imm24_20[1] ;
 wire \mod.u_cpu.cpu.immdec.imm24_20[2] ;
 wire \mod.u_cpu.cpu.immdec.imm24_20[3] ;
 wire \mod.u_cpu.cpu.immdec.imm24_20[4] ;
 wire \mod.u_cpu.cpu.immdec.imm30_25[0] ;
 wire \mod.u_cpu.cpu.immdec.imm30_25[1] ;
 wire \mod.u_cpu.cpu.immdec.imm30_25[2] ;
 wire \mod.u_cpu.cpu.immdec.imm30_25[3] ;
 wire \mod.u_cpu.cpu.immdec.imm30_25[4] ;
 wire \mod.u_cpu.cpu.immdec.imm30_25[5] ;
 wire \mod.u_cpu.cpu.immdec.imm31 ;
 wire \mod.u_cpu.cpu.immdec.imm7 ;
 wire \mod.u_cpu.cpu.mem_bytecnt[0] ;
 wire \mod.u_cpu.cpu.mem_bytecnt[1] ;
 wire \mod.u_cpu.cpu.mem_if.signbit ;
 wire \mod.u_cpu.cpu.o_wdata0 ;
 wire \mod.u_cpu.cpu.o_wdata1 ;
 wire \mod.u_cpu.cpu.o_wen0 ;
 wire \mod.u_cpu.cpu.o_wen1 ;
 wire \mod.u_cpu.cpu.state.genblk1.misalign_trap_sync_r ;
 wire \mod.u_cpu.cpu.state.ibus_cyc ;
 wire \mod.u_cpu.cpu.state.init_done ;
 wire \mod.u_cpu.cpu.state.o_cnt[2] ;
 wire \mod.u_cpu.cpu.state.o_cnt_r[0] ;
 wire \mod.u_cpu.cpu.state.o_cnt_r[1] ;
 wire \mod.u_cpu.cpu.state.o_cnt_r[2] ;
 wire \mod.u_cpu.cpu.state.o_cnt_r[3] ;
 wire \mod.u_cpu.cpu.state.stage_two_req ;
 wire \mod.u_cpu.raddr[0] ;
 wire \mod.u_cpu.raddr[1] ;
 wire \mod.u_cpu.raddr[2] ;
 wire \mod.u_cpu.raddr[3] ;
 wire \mod.u_cpu.rf_ram.memory[0][0] ;
 wire \mod.u_cpu.rf_ram.memory[0][1] ;
 wire \mod.u_cpu.rf_ram.memory[100][0] ;
 wire \mod.u_cpu.rf_ram.memory[100][1] ;
 wire \mod.u_cpu.rf_ram.memory[101][0] ;
 wire \mod.u_cpu.rf_ram.memory[101][1] ;
 wire \mod.u_cpu.rf_ram.memory[102][0] ;
 wire \mod.u_cpu.rf_ram.memory[102][1] ;
 wire \mod.u_cpu.rf_ram.memory[103][0] ;
 wire \mod.u_cpu.rf_ram.memory[103][1] ;
 wire \mod.u_cpu.rf_ram.memory[104][0] ;
 wire \mod.u_cpu.rf_ram.memory[104][1] ;
 wire \mod.u_cpu.rf_ram.memory[105][0] ;
 wire \mod.u_cpu.rf_ram.memory[105][1] ;
 wire \mod.u_cpu.rf_ram.memory[106][0] ;
 wire \mod.u_cpu.rf_ram.memory[106][1] ;
 wire \mod.u_cpu.rf_ram.memory[107][0] ;
 wire \mod.u_cpu.rf_ram.memory[107][1] ;
 wire \mod.u_cpu.rf_ram.memory[108][0] ;
 wire \mod.u_cpu.rf_ram.memory[108][1] ;
 wire \mod.u_cpu.rf_ram.memory[109][0] ;
 wire \mod.u_cpu.rf_ram.memory[109][1] ;
 wire \mod.u_cpu.rf_ram.memory[10][0] ;
 wire \mod.u_cpu.rf_ram.memory[10][1] ;
 wire \mod.u_cpu.rf_ram.memory[110][0] ;
 wire \mod.u_cpu.rf_ram.memory[110][1] ;
 wire \mod.u_cpu.rf_ram.memory[111][0] ;
 wire \mod.u_cpu.rf_ram.memory[111][1] ;
 wire \mod.u_cpu.rf_ram.memory[112][0] ;
 wire \mod.u_cpu.rf_ram.memory[112][1] ;
 wire \mod.u_cpu.rf_ram.memory[113][0] ;
 wire \mod.u_cpu.rf_ram.memory[113][1] ;
 wire \mod.u_cpu.rf_ram.memory[114][0] ;
 wire \mod.u_cpu.rf_ram.memory[114][1] ;
 wire \mod.u_cpu.rf_ram.memory[115][0] ;
 wire \mod.u_cpu.rf_ram.memory[115][1] ;
 wire \mod.u_cpu.rf_ram.memory[116][0] ;
 wire \mod.u_cpu.rf_ram.memory[116][1] ;
 wire \mod.u_cpu.rf_ram.memory[117][0] ;
 wire \mod.u_cpu.rf_ram.memory[117][1] ;
 wire \mod.u_cpu.rf_ram.memory[118][0] ;
 wire \mod.u_cpu.rf_ram.memory[118][1] ;
 wire \mod.u_cpu.rf_ram.memory[119][0] ;
 wire \mod.u_cpu.rf_ram.memory[119][1] ;
 wire \mod.u_cpu.rf_ram.memory[11][0] ;
 wire \mod.u_cpu.rf_ram.memory[11][1] ;
 wire \mod.u_cpu.rf_ram.memory[120][0] ;
 wire \mod.u_cpu.rf_ram.memory[120][1] ;
 wire \mod.u_cpu.rf_ram.memory[121][0] ;
 wire \mod.u_cpu.rf_ram.memory[121][1] ;
 wire \mod.u_cpu.rf_ram.memory[122][0] ;
 wire \mod.u_cpu.rf_ram.memory[122][1] ;
 wire \mod.u_cpu.rf_ram.memory[123][0] ;
 wire \mod.u_cpu.rf_ram.memory[123][1] ;
 wire \mod.u_cpu.rf_ram.memory[124][0] ;
 wire \mod.u_cpu.rf_ram.memory[124][1] ;
 wire \mod.u_cpu.rf_ram.memory[125][0] ;
 wire \mod.u_cpu.rf_ram.memory[125][1] ;
 wire \mod.u_cpu.rf_ram.memory[126][0] ;
 wire \mod.u_cpu.rf_ram.memory[126][1] ;
 wire \mod.u_cpu.rf_ram.memory[127][0] ;
 wire \mod.u_cpu.rf_ram.memory[127][1] ;
 wire \mod.u_cpu.rf_ram.memory[128][0] ;
 wire \mod.u_cpu.rf_ram.memory[128][1] ;
 wire \mod.u_cpu.rf_ram.memory[129][0] ;
 wire \mod.u_cpu.rf_ram.memory[129][1] ;
 wire \mod.u_cpu.rf_ram.memory[12][0] ;
 wire \mod.u_cpu.rf_ram.memory[12][1] ;
 wire \mod.u_cpu.rf_ram.memory[130][0] ;
 wire \mod.u_cpu.rf_ram.memory[130][1] ;
 wire \mod.u_cpu.rf_ram.memory[131][0] ;
 wire \mod.u_cpu.rf_ram.memory[131][1] ;
 wire \mod.u_cpu.rf_ram.memory[132][0] ;
 wire \mod.u_cpu.rf_ram.memory[132][1] ;
 wire \mod.u_cpu.rf_ram.memory[133][0] ;
 wire \mod.u_cpu.rf_ram.memory[133][1] ;
 wire \mod.u_cpu.rf_ram.memory[134][0] ;
 wire \mod.u_cpu.rf_ram.memory[134][1] ;
 wire \mod.u_cpu.rf_ram.memory[135][0] ;
 wire \mod.u_cpu.rf_ram.memory[135][1] ;
 wire \mod.u_cpu.rf_ram.memory[136][0] ;
 wire \mod.u_cpu.rf_ram.memory[136][1] ;
 wire \mod.u_cpu.rf_ram.memory[137][0] ;
 wire \mod.u_cpu.rf_ram.memory[137][1] ;
 wire \mod.u_cpu.rf_ram.memory[138][0] ;
 wire \mod.u_cpu.rf_ram.memory[138][1] ;
 wire \mod.u_cpu.rf_ram.memory[139][0] ;
 wire \mod.u_cpu.rf_ram.memory[139][1] ;
 wire \mod.u_cpu.rf_ram.memory[13][0] ;
 wire \mod.u_cpu.rf_ram.memory[13][1] ;
 wire \mod.u_cpu.rf_ram.memory[140][0] ;
 wire \mod.u_cpu.rf_ram.memory[140][1] ;
 wire \mod.u_cpu.rf_ram.memory[141][0] ;
 wire \mod.u_cpu.rf_ram.memory[141][1] ;
 wire \mod.u_cpu.rf_ram.memory[142][0] ;
 wire \mod.u_cpu.rf_ram.memory[142][1] ;
 wire \mod.u_cpu.rf_ram.memory[143][0] ;
 wire \mod.u_cpu.rf_ram.memory[143][1] ;
 wire \mod.u_cpu.rf_ram.memory[144][0] ;
 wire \mod.u_cpu.rf_ram.memory[144][1] ;
 wire \mod.u_cpu.rf_ram.memory[145][0] ;
 wire \mod.u_cpu.rf_ram.memory[145][1] ;
 wire \mod.u_cpu.rf_ram.memory[146][0] ;
 wire \mod.u_cpu.rf_ram.memory[146][1] ;
 wire \mod.u_cpu.rf_ram.memory[147][0] ;
 wire \mod.u_cpu.rf_ram.memory[147][1] ;
 wire \mod.u_cpu.rf_ram.memory[148][0] ;
 wire \mod.u_cpu.rf_ram.memory[148][1] ;
 wire \mod.u_cpu.rf_ram.memory[149][0] ;
 wire \mod.u_cpu.rf_ram.memory[149][1] ;
 wire \mod.u_cpu.rf_ram.memory[14][0] ;
 wire \mod.u_cpu.rf_ram.memory[14][1] ;
 wire \mod.u_cpu.rf_ram.memory[150][0] ;
 wire \mod.u_cpu.rf_ram.memory[150][1] ;
 wire \mod.u_cpu.rf_ram.memory[151][0] ;
 wire \mod.u_cpu.rf_ram.memory[151][1] ;
 wire \mod.u_cpu.rf_ram.memory[152][0] ;
 wire \mod.u_cpu.rf_ram.memory[152][1] ;
 wire \mod.u_cpu.rf_ram.memory[153][0] ;
 wire \mod.u_cpu.rf_ram.memory[153][1] ;
 wire \mod.u_cpu.rf_ram.memory[154][0] ;
 wire \mod.u_cpu.rf_ram.memory[154][1] ;
 wire \mod.u_cpu.rf_ram.memory[155][0] ;
 wire \mod.u_cpu.rf_ram.memory[155][1] ;
 wire \mod.u_cpu.rf_ram.memory[156][0] ;
 wire \mod.u_cpu.rf_ram.memory[156][1] ;
 wire \mod.u_cpu.rf_ram.memory[157][0] ;
 wire \mod.u_cpu.rf_ram.memory[157][1] ;
 wire \mod.u_cpu.rf_ram.memory[158][0] ;
 wire \mod.u_cpu.rf_ram.memory[158][1] ;
 wire \mod.u_cpu.rf_ram.memory[159][0] ;
 wire \mod.u_cpu.rf_ram.memory[159][1] ;
 wire \mod.u_cpu.rf_ram.memory[15][0] ;
 wire \mod.u_cpu.rf_ram.memory[15][1] ;
 wire \mod.u_cpu.rf_ram.memory[160][0] ;
 wire \mod.u_cpu.rf_ram.memory[160][1] ;
 wire \mod.u_cpu.rf_ram.memory[161][0] ;
 wire \mod.u_cpu.rf_ram.memory[161][1] ;
 wire \mod.u_cpu.rf_ram.memory[162][0] ;
 wire \mod.u_cpu.rf_ram.memory[162][1] ;
 wire \mod.u_cpu.rf_ram.memory[163][0] ;
 wire \mod.u_cpu.rf_ram.memory[163][1] ;
 wire \mod.u_cpu.rf_ram.memory[164][0] ;
 wire \mod.u_cpu.rf_ram.memory[164][1] ;
 wire \mod.u_cpu.rf_ram.memory[165][0] ;
 wire \mod.u_cpu.rf_ram.memory[165][1] ;
 wire \mod.u_cpu.rf_ram.memory[166][0] ;
 wire \mod.u_cpu.rf_ram.memory[166][1] ;
 wire \mod.u_cpu.rf_ram.memory[167][0] ;
 wire \mod.u_cpu.rf_ram.memory[167][1] ;
 wire \mod.u_cpu.rf_ram.memory[168][0] ;
 wire \mod.u_cpu.rf_ram.memory[168][1] ;
 wire \mod.u_cpu.rf_ram.memory[169][0] ;
 wire \mod.u_cpu.rf_ram.memory[169][1] ;
 wire \mod.u_cpu.rf_ram.memory[16][0] ;
 wire \mod.u_cpu.rf_ram.memory[16][1] ;
 wire \mod.u_cpu.rf_ram.memory[170][0] ;
 wire \mod.u_cpu.rf_ram.memory[170][1] ;
 wire \mod.u_cpu.rf_ram.memory[171][0] ;
 wire \mod.u_cpu.rf_ram.memory[171][1] ;
 wire \mod.u_cpu.rf_ram.memory[172][0] ;
 wire \mod.u_cpu.rf_ram.memory[172][1] ;
 wire \mod.u_cpu.rf_ram.memory[173][0] ;
 wire \mod.u_cpu.rf_ram.memory[173][1] ;
 wire \mod.u_cpu.rf_ram.memory[174][0] ;
 wire \mod.u_cpu.rf_ram.memory[174][1] ;
 wire \mod.u_cpu.rf_ram.memory[175][0] ;
 wire \mod.u_cpu.rf_ram.memory[175][1] ;
 wire \mod.u_cpu.rf_ram.memory[176][0] ;
 wire \mod.u_cpu.rf_ram.memory[176][1] ;
 wire \mod.u_cpu.rf_ram.memory[177][0] ;
 wire \mod.u_cpu.rf_ram.memory[177][1] ;
 wire \mod.u_cpu.rf_ram.memory[178][0] ;
 wire \mod.u_cpu.rf_ram.memory[178][1] ;
 wire \mod.u_cpu.rf_ram.memory[179][0] ;
 wire \mod.u_cpu.rf_ram.memory[179][1] ;
 wire \mod.u_cpu.rf_ram.memory[17][0] ;
 wire \mod.u_cpu.rf_ram.memory[17][1] ;
 wire \mod.u_cpu.rf_ram.memory[180][0] ;
 wire \mod.u_cpu.rf_ram.memory[180][1] ;
 wire \mod.u_cpu.rf_ram.memory[181][0] ;
 wire \mod.u_cpu.rf_ram.memory[181][1] ;
 wire \mod.u_cpu.rf_ram.memory[182][0] ;
 wire \mod.u_cpu.rf_ram.memory[182][1] ;
 wire \mod.u_cpu.rf_ram.memory[183][0] ;
 wire \mod.u_cpu.rf_ram.memory[183][1] ;
 wire \mod.u_cpu.rf_ram.memory[184][0] ;
 wire \mod.u_cpu.rf_ram.memory[184][1] ;
 wire \mod.u_cpu.rf_ram.memory[185][0] ;
 wire \mod.u_cpu.rf_ram.memory[185][1] ;
 wire \mod.u_cpu.rf_ram.memory[186][0] ;
 wire \mod.u_cpu.rf_ram.memory[186][1] ;
 wire \mod.u_cpu.rf_ram.memory[187][0] ;
 wire \mod.u_cpu.rf_ram.memory[187][1] ;
 wire \mod.u_cpu.rf_ram.memory[188][0] ;
 wire \mod.u_cpu.rf_ram.memory[188][1] ;
 wire \mod.u_cpu.rf_ram.memory[189][0] ;
 wire \mod.u_cpu.rf_ram.memory[189][1] ;
 wire \mod.u_cpu.rf_ram.memory[18][0] ;
 wire \mod.u_cpu.rf_ram.memory[18][1] ;
 wire \mod.u_cpu.rf_ram.memory[190][0] ;
 wire \mod.u_cpu.rf_ram.memory[190][1] ;
 wire \mod.u_cpu.rf_ram.memory[191][0] ;
 wire \mod.u_cpu.rf_ram.memory[191][1] ;
 wire \mod.u_cpu.rf_ram.memory[192][0] ;
 wire \mod.u_cpu.rf_ram.memory[192][1] ;
 wire \mod.u_cpu.rf_ram.memory[193][0] ;
 wire \mod.u_cpu.rf_ram.memory[193][1] ;
 wire \mod.u_cpu.rf_ram.memory[194][0] ;
 wire \mod.u_cpu.rf_ram.memory[194][1] ;
 wire \mod.u_cpu.rf_ram.memory[195][0] ;
 wire \mod.u_cpu.rf_ram.memory[195][1] ;
 wire \mod.u_cpu.rf_ram.memory[196][0] ;
 wire \mod.u_cpu.rf_ram.memory[196][1] ;
 wire \mod.u_cpu.rf_ram.memory[197][0] ;
 wire \mod.u_cpu.rf_ram.memory[197][1] ;
 wire \mod.u_cpu.rf_ram.memory[198][0] ;
 wire \mod.u_cpu.rf_ram.memory[198][1] ;
 wire \mod.u_cpu.rf_ram.memory[199][0] ;
 wire \mod.u_cpu.rf_ram.memory[199][1] ;
 wire \mod.u_cpu.rf_ram.memory[19][0] ;
 wire \mod.u_cpu.rf_ram.memory[19][1] ;
 wire \mod.u_cpu.rf_ram.memory[1][0] ;
 wire \mod.u_cpu.rf_ram.memory[1][1] ;
 wire \mod.u_cpu.rf_ram.memory[200][0] ;
 wire \mod.u_cpu.rf_ram.memory[200][1] ;
 wire \mod.u_cpu.rf_ram.memory[201][0] ;
 wire \mod.u_cpu.rf_ram.memory[201][1] ;
 wire \mod.u_cpu.rf_ram.memory[202][0] ;
 wire \mod.u_cpu.rf_ram.memory[202][1] ;
 wire \mod.u_cpu.rf_ram.memory[203][0] ;
 wire \mod.u_cpu.rf_ram.memory[203][1] ;
 wire \mod.u_cpu.rf_ram.memory[204][0] ;
 wire \mod.u_cpu.rf_ram.memory[204][1] ;
 wire \mod.u_cpu.rf_ram.memory[205][0] ;
 wire \mod.u_cpu.rf_ram.memory[205][1] ;
 wire \mod.u_cpu.rf_ram.memory[206][0] ;
 wire \mod.u_cpu.rf_ram.memory[206][1] ;
 wire \mod.u_cpu.rf_ram.memory[207][0] ;
 wire \mod.u_cpu.rf_ram.memory[207][1] ;
 wire \mod.u_cpu.rf_ram.memory[208][0] ;
 wire \mod.u_cpu.rf_ram.memory[208][1] ;
 wire \mod.u_cpu.rf_ram.memory[209][0] ;
 wire \mod.u_cpu.rf_ram.memory[209][1] ;
 wire \mod.u_cpu.rf_ram.memory[20][0] ;
 wire \mod.u_cpu.rf_ram.memory[20][1] ;
 wire \mod.u_cpu.rf_ram.memory[210][0] ;
 wire \mod.u_cpu.rf_ram.memory[210][1] ;
 wire \mod.u_cpu.rf_ram.memory[211][0] ;
 wire \mod.u_cpu.rf_ram.memory[211][1] ;
 wire \mod.u_cpu.rf_ram.memory[212][0] ;
 wire \mod.u_cpu.rf_ram.memory[212][1] ;
 wire \mod.u_cpu.rf_ram.memory[213][0] ;
 wire \mod.u_cpu.rf_ram.memory[213][1] ;
 wire \mod.u_cpu.rf_ram.memory[214][0] ;
 wire \mod.u_cpu.rf_ram.memory[214][1] ;
 wire \mod.u_cpu.rf_ram.memory[215][0] ;
 wire \mod.u_cpu.rf_ram.memory[215][1] ;
 wire \mod.u_cpu.rf_ram.memory[216][0] ;
 wire \mod.u_cpu.rf_ram.memory[216][1] ;
 wire \mod.u_cpu.rf_ram.memory[217][0] ;
 wire \mod.u_cpu.rf_ram.memory[217][1] ;
 wire \mod.u_cpu.rf_ram.memory[218][0] ;
 wire \mod.u_cpu.rf_ram.memory[218][1] ;
 wire \mod.u_cpu.rf_ram.memory[219][0] ;
 wire \mod.u_cpu.rf_ram.memory[219][1] ;
 wire \mod.u_cpu.rf_ram.memory[21][0] ;
 wire \mod.u_cpu.rf_ram.memory[21][1] ;
 wire \mod.u_cpu.rf_ram.memory[220][0] ;
 wire \mod.u_cpu.rf_ram.memory[220][1] ;
 wire \mod.u_cpu.rf_ram.memory[221][0] ;
 wire \mod.u_cpu.rf_ram.memory[221][1] ;
 wire \mod.u_cpu.rf_ram.memory[222][0] ;
 wire \mod.u_cpu.rf_ram.memory[222][1] ;
 wire \mod.u_cpu.rf_ram.memory[223][0] ;
 wire \mod.u_cpu.rf_ram.memory[223][1] ;
 wire \mod.u_cpu.rf_ram.memory[224][0] ;
 wire \mod.u_cpu.rf_ram.memory[224][1] ;
 wire \mod.u_cpu.rf_ram.memory[225][0] ;
 wire \mod.u_cpu.rf_ram.memory[225][1] ;
 wire \mod.u_cpu.rf_ram.memory[226][0] ;
 wire \mod.u_cpu.rf_ram.memory[226][1] ;
 wire \mod.u_cpu.rf_ram.memory[227][0] ;
 wire \mod.u_cpu.rf_ram.memory[227][1] ;
 wire \mod.u_cpu.rf_ram.memory[228][0] ;
 wire \mod.u_cpu.rf_ram.memory[228][1] ;
 wire \mod.u_cpu.rf_ram.memory[229][0] ;
 wire \mod.u_cpu.rf_ram.memory[229][1] ;
 wire \mod.u_cpu.rf_ram.memory[22][0] ;
 wire \mod.u_cpu.rf_ram.memory[22][1] ;
 wire \mod.u_cpu.rf_ram.memory[230][0] ;
 wire \mod.u_cpu.rf_ram.memory[230][1] ;
 wire \mod.u_cpu.rf_ram.memory[231][0] ;
 wire \mod.u_cpu.rf_ram.memory[231][1] ;
 wire \mod.u_cpu.rf_ram.memory[232][0] ;
 wire \mod.u_cpu.rf_ram.memory[232][1] ;
 wire \mod.u_cpu.rf_ram.memory[233][0] ;
 wire \mod.u_cpu.rf_ram.memory[233][1] ;
 wire \mod.u_cpu.rf_ram.memory[234][0] ;
 wire \mod.u_cpu.rf_ram.memory[234][1] ;
 wire \mod.u_cpu.rf_ram.memory[235][0] ;
 wire \mod.u_cpu.rf_ram.memory[235][1] ;
 wire \mod.u_cpu.rf_ram.memory[236][0] ;
 wire \mod.u_cpu.rf_ram.memory[236][1] ;
 wire \mod.u_cpu.rf_ram.memory[237][0] ;
 wire \mod.u_cpu.rf_ram.memory[237][1] ;
 wire \mod.u_cpu.rf_ram.memory[238][0] ;
 wire \mod.u_cpu.rf_ram.memory[238][1] ;
 wire \mod.u_cpu.rf_ram.memory[239][0] ;
 wire \mod.u_cpu.rf_ram.memory[239][1] ;
 wire \mod.u_cpu.rf_ram.memory[23][0] ;
 wire \mod.u_cpu.rf_ram.memory[23][1] ;
 wire \mod.u_cpu.rf_ram.memory[240][0] ;
 wire \mod.u_cpu.rf_ram.memory[240][1] ;
 wire \mod.u_cpu.rf_ram.memory[241][0] ;
 wire \mod.u_cpu.rf_ram.memory[241][1] ;
 wire \mod.u_cpu.rf_ram.memory[242][0] ;
 wire \mod.u_cpu.rf_ram.memory[242][1] ;
 wire \mod.u_cpu.rf_ram.memory[243][0] ;
 wire \mod.u_cpu.rf_ram.memory[243][1] ;
 wire \mod.u_cpu.rf_ram.memory[244][0] ;
 wire \mod.u_cpu.rf_ram.memory[244][1] ;
 wire \mod.u_cpu.rf_ram.memory[245][0] ;
 wire \mod.u_cpu.rf_ram.memory[245][1] ;
 wire \mod.u_cpu.rf_ram.memory[246][0] ;
 wire \mod.u_cpu.rf_ram.memory[246][1] ;
 wire \mod.u_cpu.rf_ram.memory[247][0] ;
 wire \mod.u_cpu.rf_ram.memory[247][1] ;
 wire \mod.u_cpu.rf_ram.memory[248][0] ;
 wire \mod.u_cpu.rf_ram.memory[248][1] ;
 wire \mod.u_cpu.rf_ram.memory[249][0] ;
 wire \mod.u_cpu.rf_ram.memory[249][1] ;
 wire \mod.u_cpu.rf_ram.memory[24][0] ;
 wire \mod.u_cpu.rf_ram.memory[24][1] ;
 wire \mod.u_cpu.rf_ram.memory[250][0] ;
 wire \mod.u_cpu.rf_ram.memory[250][1] ;
 wire \mod.u_cpu.rf_ram.memory[251][0] ;
 wire \mod.u_cpu.rf_ram.memory[251][1] ;
 wire \mod.u_cpu.rf_ram.memory[252][0] ;
 wire \mod.u_cpu.rf_ram.memory[252][1] ;
 wire \mod.u_cpu.rf_ram.memory[253][0] ;
 wire \mod.u_cpu.rf_ram.memory[253][1] ;
 wire \mod.u_cpu.rf_ram.memory[254][0] ;
 wire \mod.u_cpu.rf_ram.memory[254][1] ;
 wire \mod.u_cpu.rf_ram.memory[255][0] ;
 wire \mod.u_cpu.rf_ram.memory[255][1] ;
 wire \mod.u_cpu.rf_ram.memory[256][0] ;
 wire \mod.u_cpu.rf_ram.memory[256][1] ;
 wire \mod.u_cpu.rf_ram.memory[257][0] ;
 wire \mod.u_cpu.rf_ram.memory[257][1] ;
 wire \mod.u_cpu.rf_ram.memory[258][0] ;
 wire \mod.u_cpu.rf_ram.memory[258][1] ;
 wire \mod.u_cpu.rf_ram.memory[259][0] ;
 wire \mod.u_cpu.rf_ram.memory[259][1] ;
 wire \mod.u_cpu.rf_ram.memory[25][0] ;
 wire \mod.u_cpu.rf_ram.memory[25][1] ;
 wire \mod.u_cpu.rf_ram.memory[260][0] ;
 wire \mod.u_cpu.rf_ram.memory[260][1] ;
 wire \mod.u_cpu.rf_ram.memory[261][0] ;
 wire \mod.u_cpu.rf_ram.memory[261][1] ;
 wire \mod.u_cpu.rf_ram.memory[262][0] ;
 wire \mod.u_cpu.rf_ram.memory[262][1] ;
 wire \mod.u_cpu.rf_ram.memory[263][0] ;
 wire \mod.u_cpu.rf_ram.memory[263][1] ;
 wire \mod.u_cpu.rf_ram.memory[264][0] ;
 wire \mod.u_cpu.rf_ram.memory[264][1] ;
 wire \mod.u_cpu.rf_ram.memory[265][0] ;
 wire \mod.u_cpu.rf_ram.memory[265][1] ;
 wire \mod.u_cpu.rf_ram.memory[266][0] ;
 wire \mod.u_cpu.rf_ram.memory[266][1] ;
 wire \mod.u_cpu.rf_ram.memory[267][0] ;
 wire \mod.u_cpu.rf_ram.memory[267][1] ;
 wire \mod.u_cpu.rf_ram.memory[268][0] ;
 wire \mod.u_cpu.rf_ram.memory[268][1] ;
 wire \mod.u_cpu.rf_ram.memory[269][0] ;
 wire \mod.u_cpu.rf_ram.memory[269][1] ;
 wire \mod.u_cpu.rf_ram.memory[26][0] ;
 wire \mod.u_cpu.rf_ram.memory[26][1] ;
 wire \mod.u_cpu.rf_ram.memory[270][0] ;
 wire \mod.u_cpu.rf_ram.memory[270][1] ;
 wire \mod.u_cpu.rf_ram.memory[271][0] ;
 wire \mod.u_cpu.rf_ram.memory[271][1] ;
 wire \mod.u_cpu.rf_ram.memory[272][0] ;
 wire \mod.u_cpu.rf_ram.memory[272][1] ;
 wire \mod.u_cpu.rf_ram.memory[273][0] ;
 wire \mod.u_cpu.rf_ram.memory[273][1] ;
 wire \mod.u_cpu.rf_ram.memory[274][0] ;
 wire \mod.u_cpu.rf_ram.memory[274][1] ;
 wire \mod.u_cpu.rf_ram.memory[275][0] ;
 wire \mod.u_cpu.rf_ram.memory[275][1] ;
 wire \mod.u_cpu.rf_ram.memory[276][0] ;
 wire \mod.u_cpu.rf_ram.memory[276][1] ;
 wire \mod.u_cpu.rf_ram.memory[277][0] ;
 wire \mod.u_cpu.rf_ram.memory[277][1] ;
 wire \mod.u_cpu.rf_ram.memory[278][0] ;
 wire \mod.u_cpu.rf_ram.memory[278][1] ;
 wire \mod.u_cpu.rf_ram.memory[279][0] ;
 wire \mod.u_cpu.rf_ram.memory[279][1] ;
 wire \mod.u_cpu.rf_ram.memory[27][0] ;
 wire \mod.u_cpu.rf_ram.memory[27][1] ;
 wire \mod.u_cpu.rf_ram.memory[280][0] ;
 wire \mod.u_cpu.rf_ram.memory[280][1] ;
 wire \mod.u_cpu.rf_ram.memory[281][0] ;
 wire \mod.u_cpu.rf_ram.memory[281][1] ;
 wire \mod.u_cpu.rf_ram.memory[282][0] ;
 wire \mod.u_cpu.rf_ram.memory[282][1] ;
 wire \mod.u_cpu.rf_ram.memory[283][0] ;
 wire \mod.u_cpu.rf_ram.memory[283][1] ;
 wire \mod.u_cpu.rf_ram.memory[284][0] ;
 wire \mod.u_cpu.rf_ram.memory[284][1] ;
 wire \mod.u_cpu.rf_ram.memory[285][0] ;
 wire \mod.u_cpu.rf_ram.memory[285][1] ;
 wire \mod.u_cpu.rf_ram.memory[286][0] ;
 wire \mod.u_cpu.rf_ram.memory[286][1] ;
 wire \mod.u_cpu.rf_ram.memory[287][0] ;
 wire \mod.u_cpu.rf_ram.memory[287][1] ;
 wire \mod.u_cpu.rf_ram.memory[288][0] ;
 wire \mod.u_cpu.rf_ram.memory[288][1] ;
 wire \mod.u_cpu.rf_ram.memory[289][0] ;
 wire \mod.u_cpu.rf_ram.memory[289][1] ;
 wire \mod.u_cpu.rf_ram.memory[28][0] ;
 wire \mod.u_cpu.rf_ram.memory[28][1] ;
 wire \mod.u_cpu.rf_ram.memory[290][0] ;
 wire \mod.u_cpu.rf_ram.memory[290][1] ;
 wire \mod.u_cpu.rf_ram.memory[291][0] ;
 wire \mod.u_cpu.rf_ram.memory[291][1] ;
 wire \mod.u_cpu.rf_ram.memory[292][0] ;
 wire \mod.u_cpu.rf_ram.memory[292][1] ;
 wire \mod.u_cpu.rf_ram.memory[293][0] ;
 wire \mod.u_cpu.rf_ram.memory[293][1] ;
 wire \mod.u_cpu.rf_ram.memory[294][0] ;
 wire \mod.u_cpu.rf_ram.memory[294][1] ;
 wire \mod.u_cpu.rf_ram.memory[295][0] ;
 wire \mod.u_cpu.rf_ram.memory[295][1] ;
 wire \mod.u_cpu.rf_ram.memory[296][0] ;
 wire \mod.u_cpu.rf_ram.memory[296][1] ;
 wire \mod.u_cpu.rf_ram.memory[297][0] ;
 wire \mod.u_cpu.rf_ram.memory[297][1] ;
 wire \mod.u_cpu.rf_ram.memory[298][0] ;
 wire \mod.u_cpu.rf_ram.memory[298][1] ;
 wire \mod.u_cpu.rf_ram.memory[299][0] ;
 wire \mod.u_cpu.rf_ram.memory[299][1] ;
 wire \mod.u_cpu.rf_ram.memory[29][0] ;
 wire \mod.u_cpu.rf_ram.memory[29][1] ;
 wire \mod.u_cpu.rf_ram.memory[2][0] ;
 wire \mod.u_cpu.rf_ram.memory[2][1] ;
 wire \mod.u_cpu.rf_ram.memory[300][0] ;
 wire \mod.u_cpu.rf_ram.memory[300][1] ;
 wire \mod.u_cpu.rf_ram.memory[301][0] ;
 wire \mod.u_cpu.rf_ram.memory[301][1] ;
 wire \mod.u_cpu.rf_ram.memory[302][0] ;
 wire \mod.u_cpu.rf_ram.memory[302][1] ;
 wire \mod.u_cpu.rf_ram.memory[303][0] ;
 wire \mod.u_cpu.rf_ram.memory[303][1] ;
 wire \mod.u_cpu.rf_ram.memory[304][0] ;
 wire \mod.u_cpu.rf_ram.memory[304][1] ;
 wire \mod.u_cpu.rf_ram.memory[305][0] ;
 wire \mod.u_cpu.rf_ram.memory[305][1] ;
 wire \mod.u_cpu.rf_ram.memory[306][0] ;
 wire \mod.u_cpu.rf_ram.memory[306][1] ;
 wire \mod.u_cpu.rf_ram.memory[307][0] ;
 wire \mod.u_cpu.rf_ram.memory[307][1] ;
 wire \mod.u_cpu.rf_ram.memory[308][0] ;
 wire \mod.u_cpu.rf_ram.memory[308][1] ;
 wire \mod.u_cpu.rf_ram.memory[309][0] ;
 wire \mod.u_cpu.rf_ram.memory[309][1] ;
 wire \mod.u_cpu.rf_ram.memory[30][0] ;
 wire \mod.u_cpu.rf_ram.memory[30][1] ;
 wire \mod.u_cpu.rf_ram.memory[310][0] ;
 wire \mod.u_cpu.rf_ram.memory[310][1] ;
 wire \mod.u_cpu.rf_ram.memory[311][0] ;
 wire \mod.u_cpu.rf_ram.memory[311][1] ;
 wire \mod.u_cpu.rf_ram.memory[312][0] ;
 wire \mod.u_cpu.rf_ram.memory[312][1] ;
 wire \mod.u_cpu.rf_ram.memory[313][0] ;
 wire \mod.u_cpu.rf_ram.memory[313][1] ;
 wire \mod.u_cpu.rf_ram.memory[314][0] ;
 wire \mod.u_cpu.rf_ram.memory[314][1] ;
 wire \mod.u_cpu.rf_ram.memory[315][0] ;
 wire \mod.u_cpu.rf_ram.memory[315][1] ;
 wire \mod.u_cpu.rf_ram.memory[316][0] ;
 wire \mod.u_cpu.rf_ram.memory[316][1] ;
 wire \mod.u_cpu.rf_ram.memory[317][0] ;
 wire \mod.u_cpu.rf_ram.memory[317][1] ;
 wire \mod.u_cpu.rf_ram.memory[318][0] ;
 wire \mod.u_cpu.rf_ram.memory[318][1] ;
 wire \mod.u_cpu.rf_ram.memory[319][0] ;
 wire \mod.u_cpu.rf_ram.memory[319][1] ;
 wire \mod.u_cpu.rf_ram.memory[31][0] ;
 wire \mod.u_cpu.rf_ram.memory[31][1] ;
 wire \mod.u_cpu.rf_ram.memory[320][0] ;
 wire \mod.u_cpu.rf_ram.memory[320][1] ;
 wire \mod.u_cpu.rf_ram.memory[321][0] ;
 wire \mod.u_cpu.rf_ram.memory[321][1] ;
 wire \mod.u_cpu.rf_ram.memory[322][0] ;
 wire \mod.u_cpu.rf_ram.memory[322][1] ;
 wire \mod.u_cpu.rf_ram.memory[323][0] ;
 wire \mod.u_cpu.rf_ram.memory[323][1] ;
 wire \mod.u_cpu.rf_ram.memory[324][0] ;
 wire \mod.u_cpu.rf_ram.memory[324][1] ;
 wire \mod.u_cpu.rf_ram.memory[325][0] ;
 wire \mod.u_cpu.rf_ram.memory[325][1] ;
 wire \mod.u_cpu.rf_ram.memory[326][0] ;
 wire \mod.u_cpu.rf_ram.memory[326][1] ;
 wire \mod.u_cpu.rf_ram.memory[327][0] ;
 wire \mod.u_cpu.rf_ram.memory[327][1] ;
 wire \mod.u_cpu.rf_ram.memory[328][0] ;
 wire \mod.u_cpu.rf_ram.memory[328][1] ;
 wire \mod.u_cpu.rf_ram.memory[329][0] ;
 wire \mod.u_cpu.rf_ram.memory[329][1] ;
 wire \mod.u_cpu.rf_ram.memory[32][0] ;
 wire \mod.u_cpu.rf_ram.memory[32][1] ;
 wire \mod.u_cpu.rf_ram.memory[330][0] ;
 wire \mod.u_cpu.rf_ram.memory[330][1] ;
 wire \mod.u_cpu.rf_ram.memory[331][0] ;
 wire \mod.u_cpu.rf_ram.memory[331][1] ;
 wire \mod.u_cpu.rf_ram.memory[332][0] ;
 wire \mod.u_cpu.rf_ram.memory[332][1] ;
 wire \mod.u_cpu.rf_ram.memory[333][0] ;
 wire \mod.u_cpu.rf_ram.memory[333][1] ;
 wire \mod.u_cpu.rf_ram.memory[334][0] ;
 wire \mod.u_cpu.rf_ram.memory[334][1] ;
 wire \mod.u_cpu.rf_ram.memory[335][0] ;
 wire \mod.u_cpu.rf_ram.memory[335][1] ;
 wire \mod.u_cpu.rf_ram.memory[336][0] ;
 wire \mod.u_cpu.rf_ram.memory[336][1] ;
 wire \mod.u_cpu.rf_ram.memory[337][0] ;
 wire \mod.u_cpu.rf_ram.memory[337][1] ;
 wire \mod.u_cpu.rf_ram.memory[338][0] ;
 wire \mod.u_cpu.rf_ram.memory[338][1] ;
 wire \mod.u_cpu.rf_ram.memory[339][0] ;
 wire \mod.u_cpu.rf_ram.memory[339][1] ;
 wire \mod.u_cpu.rf_ram.memory[33][0] ;
 wire \mod.u_cpu.rf_ram.memory[33][1] ;
 wire \mod.u_cpu.rf_ram.memory[340][0] ;
 wire \mod.u_cpu.rf_ram.memory[340][1] ;
 wire \mod.u_cpu.rf_ram.memory[341][0] ;
 wire \mod.u_cpu.rf_ram.memory[341][1] ;
 wire \mod.u_cpu.rf_ram.memory[342][0] ;
 wire \mod.u_cpu.rf_ram.memory[342][1] ;
 wire \mod.u_cpu.rf_ram.memory[343][0] ;
 wire \mod.u_cpu.rf_ram.memory[343][1] ;
 wire \mod.u_cpu.rf_ram.memory[344][0] ;
 wire \mod.u_cpu.rf_ram.memory[344][1] ;
 wire \mod.u_cpu.rf_ram.memory[345][0] ;
 wire \mod.u_cpu.rf_ram.memory[345][1] ;
 wire \mod.u_cpu.rf_ram.memory[346][0] ;
 wire \mod.u_cpu.rf_ram.memory[346][1] ;
 wire \mod.u_cpu.rf_ram.memory[347][0] ;
 wire \mod.u_cpu.rf_ram.memory[347][1] ;
 wire \mod.u_cpu.rf_ram.memory[348][0] ;
 wire \mod.u_cpu.rf_ram.memory[348][1] ;
 wire \mod.u_cpu.rf_ram.memory[349][0] ;
 wire \mod.u_cpu.rf_ram.memory[349][1] ;
 wire \mod.u_cpu.rf_ram.memory[34][0] ;
 wire \mod.u_cpu.rf_ram.memory[34][1] ;
 wire \mod.u_cpu.rf_ram.memory[350][0] ;
 wire \mod.u_cpu.rf_ram.memory[350][1] ;
 wire \mod.u_cpu.rf_ram.memory[351][0] ;
 wire \mod.u_cpu.rf_ram.memory[351][1] ;
 wire \mod.u_cpu.rf_ram.memory[352][0] ;
 wire \mod.u_cpu.rf_ram.memory[352][1] ;
 wire \mod.u_cpu.rf_ram.memory[353][0] ;
 wire \mod.u_cpu.rf_ram.memory[353][1] ;
 wire \mod.u_cpu.rf_ram.memory[354][0] ;
 wire \mod.u_cpu.rf_ram.memory[354][1] ;
 wire \mod.u_cpu.rf_ram.memory[355][0] ;
 wire \mod.u_cpu.rf_ram.memory[355][1] ;
 wire \mod.u_cpu.rf_ram.memory[356][0] ;
 wire \mod.u_cpu.rf_ram.memory[356][1] ;
 wire \mod.u_cpu.rf_ram.memory[357][0] ;
 wire \mod.u_cpu.rf_ram.memory[357][1] ;
 wire \mod.u_cpu.rf_ram.memory[358][0] ;
 wire \mod.u_cpu.rf_ram.memory[358][1] ;
 wire \mod.u_cpu.rf_ram.memory[359][0] ;
 wire \mod.u_cpu.rf_ram.memory[359][1] ;
 wire \mod.u_cpu.rf_ram.memory[35][0] ;
 wire \mod.u_cpu.rf_ram.memory[35][1] ;
 wire \mod.u_cpu.rf_ram.memory[360][0] ;
 wire \mod.u_cpu.rf_ram.memory[360][1] ;
 wire \mod.u_cpu.rf_ram.memory[361][0] ;
 wire \mod.u_cpu.rf_ram.memory[361][1] ;
 wire \mod.u_cpu.rf_ram.memory[362][0] ;
 wire \mod.u_cpu.rf_ram.memory[362][1] ;
 wire \mod.u_cpu.rf_ram.memory[363][0] ;
 wire \mod.u_cpu.rf_ram.memory[363][1] ;
 wire \mod.u_cpu.rf_ram.memory[364][0] ;
 wire \mod.u_cpu.rf_ram.memory[364][1] ;
 wire \mod.u_cpu.rf_ram.memory[365][0] ;
 wire \mod.u_cpu.rf_ram.memory[365][1] ;
 wire \mod.u_cpu.rf_ram.memory[366][0] ;
 wire \mod.u_cpu.rf_ram.memory[366][1] ;
 wire \mod.u_cpu.rf_ram.memory[367][0] ;
 wire \mod.u_cpu.rf_ram.memory[367][1] ;
 wire \mod.u_cpu.rf_ram.memory[368][0] ;
 wire \mod.u_cpu.rf_ram.memory[368][1] ;
 wire \mod.u_cpu.rf_ram.memory[369][0] ;
 wire \mod.u_cpu.rf_ram.memory[369][1] ;
 wire \mod.u_cpu.rf_ram.memory[36][0] ;
 wire \mod.u_cpu.rf_ram.memory[36][1] ;
 wire \mod.u_cpu.rf_ram.memory[370][0] ;
 wire \mod.u_cpu.rf_ram.memory[370][1] ;
 wire \mod.u_cpu.rf_ram.memory[371][0] ;
 wire \mod.u_cpu.rf_ram.memory[371][1] ;
 wire \mod.u_cpu.rf_ram.memory[372][0] ;
 wire \mod.u_cpu.rf_ram.memory[372][1] ;
 wire \mod.u_cpu.rf_ram.memory[373][0] ;
 wire \mod.u_cpu.rf_ram.memory[373][1] ;
 wire \mod.u_cpu.rf_ram.memory[374][0] ;
 wire \mod.u_cpu.rf_ram.memory[374][1] ;
 wire \mod.u_cpu.rf_ram.memory[375][0] ;
 wire \mod.u_cpu.rf_ram.memory[375][1] ;
 wire \mod.u_cpu.rf_ram.memory[376][0] ;
 wire \mod.u_cpu.rf_ram.memory[376][1] ;
 wire \mod.u_cpu.rf_ram.memory[377][0] ;
 wire \mod.u_cpu.rf_ram.memory[377][1] ;
 wire \mod.u_cpu.rf_ram.memory[378][0] ;
 wire \mod.u_cpu.rf_ram.memory[378][1] ;
 wire \mod.u_cpu.rf_ram.memory[379][0] ;
 wire \mod.u_cpu.rf_ram.memory[379][1] ;
 wire \mod.u_cpu.rf_ram.memory[37][0] ;
 wire \mod.u_cpu.rf_ram.memory[37][1] ;
 wire \mod.u_cpu.rf_ram.memory[380][0] ;
 wire \mod.u_cpu.rf_ram.memory[380][1] ;
 wire \mod.u_cpu.rf_ram.memory[381][0] ;
 wire \mod.u_cpu.rf_ram.memory[381][1] ;
 wire \mod.u_cpu.rf_ram.memory[382][0] ;
 wire \mod.u_cpu.rf_ram.memory[382][1] ;
 wire \mod.u_cpu.rf_ram.memory[383][0] ;
 wire \mod.u_cpu.rf_ram.memory[383][1] ;
 wire \mod.u_cpu.rf_ram.memory[384][0] ;
 wire \mod.u_cpu.rf_ram.memory[384][1] ;
 wire \mod.u_cpu.rf_ram.memory[385][0] ;
 wire \mod.u_cpu.rf_ram.memory[385][1] ;
 wire \mod.u_cpu.rf_ram.memory[386][0] ;
 wire \mod.u_cpu.rf_ram.memory[386][1] ;
 wire \mod.u_cpu.rf_ram.memory[387][0] ;
 wire \mod.u_cpu.rf_ram.memory[387][1] ;
 wire \mod.u_cpu.rf_ram.memory[388][0] ;
 wire \mod.u_cpu.rf_ram.memory[388][1] ;
 wire \mod.u_cpu.rf_ram.memory[389][0] ;
 wire \mod.u_cpu.rf_ram.memory[389][1] ;
 wire \mod.u_cpu.rf_ram.memory[38][0] ;
 wire \mod.u_cpu.rf_ram.memory[38][1] ;
 wire \mod.u_cpu.rf_ram.memory[390][0] ;
 wire \mod.u_cpu.rf_ram.memory[390][1] ;
 wire \mod.u_cpu.rf_ram.memory[391][0] ;
 wire \mod.u_cpu.rf_ram.memory[391][1] ;
 wire \mod.u_cpu.rf_ram.memory[392][0] ;
 wire \mod.u_cpu.rf_ram.memory[392][1] ;
 wire \mod.u_cpu.rf_ram.memory[393][0] ;
 wire \mod.u_cpu.rf_ram.memory[393][1] ;
 wire \mod.u_cpu.rf_ram.memory[394][0] ;
 wire \mod.u_cpu.rf_ram.memory[394][1] ;
 wire \mod.u_cpu.rf_ram.memory[395][0] ;
 wire \mod.u_cpu.rf_ram.memory[395][1] ;
 wire \mod.u_cpu.rf_ram.memory[396][0] ;
 wire \mod.u_cpu.rf_ram.memory[396][1] ;
 wire \mod.u_cpu.rf_ram.memory[397][0] ;
 wire \mod.u_cpu.rf_ram.memory[397][1] ;
 wire \mod.u_cpu.rf_ram.memory[398][0] ;
 wire \mod.u_cpu.rf_ram.memory[398][1] ;
 wire \mod.u_cpu.rf_ram.memory[399][0] ;
 wire \mod.u_cpu.rf_ram.memory[399][1] ;
 wire \mod.u_cpu.rf_ram.memory[39][0] ;
 wire \mod.u_cpu.rf_ram.memory[39][1] ;
 wire \mod.u_cpu.rf_ram.memory[3][0] ;
 wire \mod.u_cpu.rf_ram.memory[3][1] ;
 wire \mod.u_cpu.rf_ram.memory[400][0] ;
 wire \mod.u_cpu.rf_ram.memory[400][1] ;
 wire \mod.u_cpu.rf_ram.memory[401][0] ;
 wire \mod.u_cpu.rf_ram.memory[401][1] ;
 wire \mod.u_cpu.rf_ram.memory[402][0] ;
 wire \mod.u_cpu.rf_ram.memory[402][1] ;
 wire \mod.u_cpu.rf_ram.memory[403][0] ;
 wire \mod.u_cpu.rf_ram.memory[403][1] ;
 wire \mod.u_cpu.rf_ram.memory[404][0] ;
 wire \mod.u_cpu.rf_ram.memory[404][1] ;
 wire \mod.u_cpu.rf_ram.memory[405][0] ;
 wire \mod.u_cpu.rf_ram.memory[405][1] ;
 wire \mod.u_cpu.rf_ram.memory[406][0] ;
 wire \mod.u_cpu.rf_ram.memory[406][1] ;
 wire \mod.u_cpu.rf_ram.memory[407][0] ;
 wire \mod.u_cpu.rf_ram.memory[407][1] ;
 wire \mod.u_cpu.rf_ram.memory[408][0] ;
 wire \mod.u_cpu.rf_ram.memory[408][1] ;
 wire \mod.u_cpu.rf_ram.memory[409][0] ;
 wire \mod.u_cpu.rf_ram.memory[409][1] ;
 wire \mod.u_cpu.rf_ram.memory[40][0] ;
 wire \mod.u_cpu.rf_ram.memory[40][1] ;
 wire \mod.u_cpu.rf_ram.memory[410][0] ;
 wire \mod.u_cpu.rf_ram.memory[410][1] ;
 wire \mod.u_cpu.rf_ram.memory[411][0] ;
 wire \mod.u_cpu.rf_ram.memory[411][1] ;
 wire \mod.u_cpu.rf_ram.memory[412][0] ;
 wire \mod.u_cpu.rf_ram.memory[412][1] ;
 wire \mod.u_cpu.rf_ram.memory[413][0] ;
 wire \mod.u_cpu.rf_ram.memory[413][1] ;
 wire \mod.u_cpu.rf_ram.memory[414][0] ;
 wire \mod.u_cpu.rf_ram.memory[414][1] ;
 wire \mod.u_cpu.rf_ram.memory[415][0] ;
 wire \mod.u_cpu.rf_ram.memory[415][1] ;
 wire \mod.u_cpu.rf_ram.memory[416][0] ;
 wire \mod.u_cpu.rf_ram.memory[416][1] ;
 wire \mod.u_cpu.rf_ram.memory[417][0] ;
 wire \mod.u_cpu.rf_ram.memory[417][1] ;
 wire \mod.u_cpu.rf_ram.memory[418][0] ;
 wire \mod.u_cpu.rf_ram.memory[418][1] ;
 wire \mod.u_cpu.rf_ram.memory[419][0] ;
 wire \mod.u_cpu.rf_ram.memory[419][1] ;
 wire \mod.u_cpu.rf_ram.memory[41][0] ;
 wire \mod.u_cpu.rf_ram.memory[41][1] ;
 wire \mod.u_cpu.rf_ram.memory[420][0] ;
 wire \mod.u_cpu.rf_ram.memory[420][1] ;
 wire \mod.u_cpu.rf_ram.memory[421][0] ;
 wire \mod.u_cpu.rf_ram.memory[421][1] ;
 wire \mod.u_cpu.rf_ram.memory[422][0] ;
 wire \mod.u_cpu.rf_ram.memory[422][1] ;
 wire \mod.u_cpu.rf_ram.memory[423][0] ;
 wire \mod.u_cpu.rf_ram.memory[423][1] ;
 wire \mod.u_cpu.rf_ram.memory[424][0] ;
 wire \mod.u_cpu.rf_ram.memory[424][1] ;
 wire \mod.u_cpu.rf_ram.memory[425][0] ;
 wire \mod.u_cpu.rf_ram.memory[425][1] ;
 wire \mod.u_cpu.rf_ram.memory[426][0] ;
 wire \mod.u_cpu.rf_ram.memory[426][1] ;
 wire \mod.u_cpu.rf_ram.memory[427][0] ;
 wire \mod.u_cpu.rf_ram.memory[427][1] ;
 wire \mod.u_cpu.rf_ram.memory[428][0] ;
 wire \mod.u_cpu.rf_ram.memory[428][1] ;
 wire \mod.u_cpu.rf_ram.memory[429][0] ;
 wire \mod.u_cpu.rf_ram.memory[429][1] ;
 wire \mod.u_cpu.rf_ram.memory[42][0] ;
 wire \mod.u_cpu.rf_ram.memory[42][1] ;
 wire \mod.u_cpu.rf_ram.memory[430][0] ;
 wire \mod.u_cpu.rf_ram.memory[430][1] ;
 wire \mod.u_cpu.rf_ram.memory[431][0] ;
 wire \mod.u_cpu.rf_ram.memory[431][1] ;
 wire \mod.u_cpu.rf_ram.memory[432][0] ;
 wire \mod.u_cpu.rf_ram.memory[432][1] ;
 wire \mod.u_cpu.rf_ram.memory[433][0] ;
 wire \mod.u_cpu.rf_ram.memory[433][1] ;
 wire \mod.u_cpu.rf_ram.memory[434][0] ;
 wire \mod.u_cpu.rf_ram.memory[434][1] ;
 wire \mod.u_cpu.rf_ram.memory[435][0] ;
 wire \mod.u_cpu.rf_ram.memory[435][1] ;
 wire \mod.u_cpu.rf_ram.memory[436][0] ;
 wire \mod.u_cpu.rf_ram.memory[436][1] ;
 wire \mod.u_cpu.rf_ram.memory[437][0] ;
 wire \mod.u_cpu.rf_ram.memory[437][1] ;
 wire \mod.u_cpu.rf_ram.memory[438][0] ;
 wire \mod.u_cpu.rf_ram.memory[438][1] ;
 wire \mod.u_cpu.rf_ram.memory[439][0] ;
 wire \mod.u_cpu.rf_ram.memory[439][1] ;
 wire \mod.u_cpu.rf_ram.memory[43][0] ;
 wire \mod.u_cpu.rf_ram.memory[43][1] ;
 wire \mod.u_cpu.rf_ram.memory[440][0] ;
 wire \mod.u_cpu.rf_ram.memory[440][1] ;
 wire \mod.u_cpu.rf_ram.memory[441][0] ;
 wire \mod.u_cpu.rf_ram.memory[441][1] ;
 wire \mod.u_cpu.rf_ram.memory[442][0] ;
 wire \mod.u_cpu.rf_ram.memory[442][1] ;
 wire \mod.u_cpu.rf_ram.memory[443][0] ;
 wire \mod.u_cpu.rf_ram.memory[443][1] ;
 wire \mod.u_cpu.rf_ram.memory[444][0] ;
 wire \mod.u_cpu.rf_ram.memory[444][1] ;
 wire \mod.u_cpu.rf_ram.memory[445][0] ;
 wire \mod.u_cpu.rf_ram.memory[445][1] ;
 wire \mod.u_cpu.rf_ram.memory[446][0] ;
 wire \mod.u_cpu.rf_ram.memory[446][1] ;
 wire \mod.u_cpu.rf_ram.memory[447][0] ;
 wire \mod.u_cpu.rf_ram.memory[447][1] ;
 wire \mod.u_cpu.rf_ram.memory[448][0] ;
 wire \mod.u_cpu.rf_ram.memory[448][1] ;
 wire \mod.u_cpu.rf_ram.memory[449][0] ;
 wire \mod.u_cpu.rf_ram.memory[449][1] ;
 wire \mod.u_cpu.rf_ram.memory[44][0] ;
 wire \mod.u_cpu.rf_ram.memory[44][1] ;
 wire \mod.u_cpu.rf_ram.memory[450][0] ;
 wire \mod.u_cpu.rf_ram.memory[450][1] ;
 wire \mod.u_cpu.rf_ram.memory[451][0] ;
 wire \mod.u_cpu.rf_ram.memory[451][1] ;
 wire \mod.u_cpu.rf_ram.memory[452][0] ;
 wire \mod.u_cpu.rf_ram.memory[452][1] ;
 wire \mod.u_cpu.rf_ram.memory[453][0] ;
 wire \mod.u_cpu.rf_ram.memory[453][1] ;
 wire \mod.u_cpu.rf_ram.memory[454][0] ;
 wire \mod.u_cpu.rf_ram.memory[454][1] ;
 wire \mod.u_cpu.rf_ram.memory[455][0] ;
 wire \mod.u_cpu.rf_ram.memory[455][1] ;
 wire \mod.u_cpu.rf_ram.memory[456][0] ;
 wire \mod.u_cpu.rf_ram.memory[456][1] ;
 wire \mod.u_cpu.rf_ram.memory[457][0] ;
 wire \mod.u_cpu.rf_ram.memory[457][1] ;
 wire \mod.u_cpu.rf_ram.memory[458][0] ;
 wire \mod.u_cpu.rf_ram.memory[458][1] ;
 wire \mod.u_cpu.rf_ram.memory[459][0] ;
 wire \mod.u_cpu.rf_ram.memory[459][1] ;
 wire \mod.u_cpu.rf_ram.memory[45][0] ;
 wire \mod.u_cpu.rf_ram.memory[45][1] ;
 wire \mod.u_cpu.rf_ram.memory[460][0] ;
 wire \mod.u_cpu.rf_ram.memory[460][1] ;
 wire \mod.u_cpu.rf_ram.memory[461][0] ;
 wire \mod.u_cpu.rf_ram.memory[461][1] ;
 wire \mod.u_cpu.rf_ram.memory[462][0] ;
 wire \mod.u_cpu.rf_ram.memory[462][1] ;
 wire \mod.u_cpu.rf_ram.memory[463][0] ;
 wire \mod.u_cpu.rf_ram.memory[463][1] ;
 wire \mod.u_cpu.rf_ram.memory[464][0] ;
 wire \mod.u_cpu.rf_ram.memory[464][1] ;
 wire \mod.u_cpu.rf_ram.memory[465][0] ;
 wire \mod.u_cpu.rf_ram.memory[465][1] ;
 wire \mod.u_cpu.rf_ram.memory[466][0] ;
 wire \mod.u_cpu.rf_ram.memory[466][1] ;
 wire \mod.u_cpu.rf_ram.memory[467][0] ;
 wire \mod.u_cpu.rf_ram.memory[467][1] ;
 wire \mod.u_cpu.rf_ram.memory[468][0] ;
 wire \mod.u_cpu.rf_ram.memory[468][1] ;
 wire \mod.u_cpu.rf_ram.memory[469][0] ;
 wire \mod.u_cpu.rf_ram.memory[469][1] ;
 wire \mod.u_cpu.rf_ram.memory[46][0] ;
 wire \mod.u_cpu.rf_ram.memory[46][1] ;
 wire \mod.u_cpu.rf_ram.memory[470][0] ;
 wire \mod.u_cpu.rf_ram.memory[470][1] ;
 wire \mod.u_cpu.rf_ram.memory[471][0] ;
 wire \mod.u_cpu.rf_ram.memory[471][1] ;
 wire \mod.u_cpu.rf_ram.memory[472][0] ;
 wire \mod.u_cpu.rf_ram.memory[472][1] ;
 wire \mod.u_cpu.rf_ram.memory[473][0] ;
 wire \mod.u_cpu.rf_ram.memory[473][1] ;
 wire \mod.u_cpu.rf_ram.memory[474][0] ;
 wire \mod.u_cpu.rf_ram.memory[474][1] ;
 wire \mod.u_cpu.rf_ram.memory[475][0] ;
 wire \mod.u_cpu.rf_ram.memory[475][1] ;
 wire \mod.u_cpu.rf_ram.memory[476][0] ;
 wire \mod.u_cpu.rf_ram.memory[476][1] ;
 wire \mod.u_cpu.rf_ram.memory[477][0] ;
 wire \mod.u_cpu.rf_ram.memory[477][1] ;
 wire \mod.u_cpu.rf_ram.memory[478][0] ;
 wire \mod.u_cpu.rf_ram.memory[478][1] ;
 wire \mod.u_cpu.rf_ram.memory[479][0] ;
 wire \mod.u_cpu.rf_ram.memory[479][1] ;
 wire \mod.u_cpu.rf_ram.memory[47][0] ;
 wire \mod.u_cpu.rf_ram.memory[47][1] ;
 wire \mod.u_cpu.rf_ram.memory[480][0] ;
 wire \mod.u_cpu.rf_ram.memory[480][1] ;
 wire \mod.u_cpu.rf_ram.memory[481][0] ;
 wire \mod.u_cpu.rf_ram.memory[481][1] ;
 wire \mod.u_cpu.rf_ram.memory[482][0] ;
 wire \mod.u_cpu.rf_ram.memory[482][1] ;
 wire \mod.u_cpu.rf_ram.memory[483][0] ;
 wire \mod.u_cpu.rf_ram.memory[483][1] ;
 wire \mod.u_cpu.rf_ram.memory[484][0] ;
 wire \mod.u_cpu.rf_ram.memory[484][1] ;
 wire \mod.u_cpu.rf_ram.memory[485][0] ;
 wire \mod.u_cpu.rf_ram.memory[485][1] ;
 wire \mod.u_cpu.rf_ram.memory[486][0] ;
 wire \mod.u_cpu.rf_ram.memory[486][1] ;
 wire \mod.u_cpu.rf_ram.memory[487][0] ;
 wire \mod.u_cpu.rf_ram.memory[487][1] ;
 wire \mod.u_cpu.rf_ram.memory[488][0] ;
 wire \mod.u_cpu.rf_ram.memory[488][1] ;
 wire \mod.u_cpu.rf_ram.memory[489][0] ;
 wire \mod.u_cpu.rf_ram.memory[489][1] ;
 wire \mod.u_cpu.rf_ram.memory[48][0] ;
 wire \mod.u_cpu.rf_ram.memory[48][1] ;
 wire \mod.u_cpu.rf_ram.memory[490][0] ;
 wire \mod.u_cpu.rf_ram.memory[490][1] ;
 wire \mod.u_cpu.rf_ram.memory[491][0] ;
 wire \mod.u_cpu.rf_ram.memory[491][1] ;
 wire \mod.u_cpu.rf_ram.memory[492][0] ;
 wire \mod.u_cpu.rf_ram.memory[492][1] ;
 wire \mod.u_cpu.rf_ram.memory[493][0] ;
 wire \mod.u_cpu.rf_ram.memory[493][1] ;
 wire \mod.u_cpu.rf_ram.memory[494][0] ;
 wire \mod.u_cpu.rf_ram.memory[494][1] ;
 wire \mod.u_cpu.rf_ram.memory[495][0] ;
 wire \mod.u_cpu.rf_ram.memory[495][1] ;
 wire \mod.u_cpu.rf_ram.memory[496][0] ;
 wire \mod.u_cpu.rf_ram.memory[496][1] ;
 wire \mod.u_cpu.rf_ram.memory[497][0] ;
 wire \mod.u_cpu.rf_ram.memory[497][1] ;
 wire \mod.u_cpu.rf_ram.memory[498][0] ;
 wire \mod.u_cpu.rf_ram.memory[498][1] ;
 wire \mod.u_cpu.rf_ram.memory[499][0] ;
 wire \mod.u_cpu.rf_ram.memory[499][1] ;
 wire \mod.u_cpu.rf_ram.memory[49][0] ;
 wire \mod.u_cpu.rf_ram.memory[49][1] ;
 wire \mod.u_cpu.rf_ram.memory[4][0] ;
 wire \mod.u_cpu.rf_ram.memory[4][1] ;
 wire \mod.u_cpu.rf_ram.memory[500][0] ;
 wire \mod.u_cpu.rf_ram.memory[500][1] ;
 wire \mod.u_cpu.rf_ram.memory[501][0] ;
 wire \mod.u_cpu.rf_ram.memory[501][1] ;
 wire \mod.u_cpu.rf_ram.memory[502][0] ;
 wire \mod.u_cpu.rf_ram.memory[502][1] ;
 wire \mod.u_cpu.rf_ram.memory[503][0] ;
 wire \mod.u_cpu.rf_ram.memory[503][1] ;
 wire \mod.u_cpu.rf_ram.memory[504][0] ;
 wire \mod.u_cpu.rf_ram.memory[504][1] ;
 wire \mod.u_cpu.rf_ram.memory[505][0] ;
 wire \mod.u_cpu.rf_ram.memory[505][1] ;
 wire \mod.u_cpu.rf_ram.memory[506][0] ;
 wire \mod.u_cpu.rf_ram.memory[506][1] ;
 wire \mod.u_cpu.rf_ram.memory[507][0] ;
 wire \mod.u_cpu.rf_ram.memory[507][1] ;
 wire \mod.u_cpu.rf_ram.memory[508][0] ;
 wire \mod.u_cpu.rf_ram.memory[508][1] ;
 wire \mod.u_cpu.rf_ram.memory[509][0] ;
 wire \mod.u_cpu.rf_ram.memory[509][1] ;
 wire \mod.u_cpu.rf_ram.memory[50][0] ;
 wire \mod.u_cpu.rf_ram.memory[50][1] ;
 wire \mod.u_cpu.rf_ram.memory[510][0] ;
 wire \mod.u_cpu.rf_ram.memory[510][1] ;
 wire \mod.u_cpu.rf_ram.memory[511][0] ;
 wire \mod.u_cpu.rf_ram.memory[511][1] ;
 wire \mod.u_cpu.rf_ram.memory[512][0] ;
 wire \mod.u_cpu.rf_ram.memory[512][1] ;
 wire \mod.u_cpu.rf_ram.memory[513][0] ;
 wire \mod.u_cpu.rf_ram.memory[513][1] ;
 wire \mod.u_cpu.rf_ram.memory[514][0] ;
 wire \mod.u_cpu.rf_ram.memory[514][1] ;
 wire \mod.u_cpu.rf_ram.memory[515][0] ;
 wire \mod.u_cpu.rf_ram.memory[515][1] ;
 wire \mod.u_cpu.rf_ram.memory[516][0] ;
 wire \mod.u_cpu.rf_ram.memory[516][1] ;
 wire \mod.u_cpu.rf_ram.memory[517][0] ;
 wire \mod.u_cpu.rf_ram.memory[517][1] ;
 wire \mod.u_cpu.rf_ram.memory[518][0] ;
 wire \mod.u_cpu.rf_ram.memory[518][1] ;
 wire \mod.u_cpu.rf_ram.memory[519][0] ;
 wire \mod.u_cpu.rf_ram.memory[519][1] ;
 wire \mod.u_cpu.rf_ram.memory[51][0] ;
 wire \mod.u_cpu.rf_ram.memory[51][1] ;
 wire \mod.u_cpu.rf_ram.memory[520][0] ;
 wire \mod.u_cpu.rf_ram.memory[520][1] ;
 wire \mod.u_cpu.rf_ram.memory[521][0] ;
 wire \mod.u_cpu.rf_ram.memory[521][1] ;
 wire \mod.u_cpu.rf_ram.memory[522][0] ;
 wire \mod.u_cpu.rf_ram.memory[522][1] ;
 wire \mod.u_cpu.rf_ram.memory[523][0] ;
 wire \mod.u_cpu.rf_ram.memory[523][1] ;
 wire \mod.u_cpu.rf_ram.memory[524][0] ;
 wire \mod.u_cpu.rf_ram.memory[524][1] ;
 wire \mod.u_cpu.rf_ram.memory[525][0] ;
 wire \mod.u_cpu.rf_ram.memory[525][1] ;
 wire \mod.u_cpu.rf_ram.memory[526][0] ;
 wire \mod.u_cpu.rf_ram.memory[526][1] ;
 wire \mod.u_cpu.rf_ram.memory[527][0] ;
 wire \mod.u_cpu.rf_ram.memory[527][1] ;
 wire \mod.u_cpu.rf_ram.memory[528][0] ;
 wire \mod.u_cpu.rf_ram.memory[528][1] ;
 wire \mod.u_cpu.rf_ram.memory[529][0] ;
 wire \mod.u_cpu.rf_ram.memory[529][1] ;
 wire \mod.u_cpu.rf_ram.memory[52][0] ;
 wire \mod.u_cpu.rf_ram.memory[52][1] ;
 wire \mod.u_cpu.rf_ram.memory[530][0] ;
 wire \mod.u_cpu.rf_ram.memory[530][1] ;
 wire \mod.u_cpu.rf_ram.memory[531][0] ;
 wire \mod.u_cpu.rf_ram.memory[531][1] ;
 wire \mod.u_cpu.rf_ram.memory[532][0] ;
 wire \mod.u_cpu.rf_ram.memory[532][1] ;
 wire \mod.u_cpu.rf_ram.memory[533][0] ;
 wire \mod.u_cpu.rf_ram.memory[533][1] ;
 wire \mod.u_cpu.rf_ram.memory[534][0] ;
 wire \mod.u_cpu.rf_ram.memory[534][1] ;
 wire \mod.u_cpu.rf_ram.memory[535][0] ;
 wire \mod.u_cpu.rf_ram.memory[535][1] ;
 wire \mod.u_cpu.rf_ram.memory[536][0] ;
 wire \mod.u_cpu.rf_ram.memory[536][1] ;
 wire \mod.u_cpu.rf_ram.memory[537][0] ;
 wire \mod.u_cpu.rf_ram.memory[537][1] ;
 wire \mod.u_cpu.rf_ram.memory[538][0] ;
 wire \mod.u_cpu.rf_ram.memory[538][1] ;
 wire \mod.u_cpu.rf_ram.memory[539][0] ;
 wire \mod.u_cpu.rf_ram.memory[539][1] ;
 wire \mod.u_cpu.rf_ram.memory[53][0] ;
 wire \mod.u_cpu.rf_ram.memory[53][1] ;
 wire \mod.u_cpu.rf_ram.memory[540][0] ;
 wire \mod.u_cpu.rf_ram.memory[540][1] ;
 wire \mod.u_cpu.rf_ram.memory[541][0] ;
 wire \mod.u_cpu.rf_ram.memory[541][1] ;
 wire \mod.u_cpu.rf_ram.memory[542][0] ;
 wire \mod.u_cpu.rf_ram.memory[542][1] ;
 wire \mod.u_cpu.rf_ram.memory[543][0] ;
 wire \mod.u_cpu.rf_ram.memory[543][1] ;
 wire \mod.u_cpu.rf_ram.memory[544][0] ;
 wire \mod.u_cpu.rf_ram.memory[544][1] ;
 wire \mod.u_cpu.rf_ram.memory[545][0] ;
 wire \mod.u_cpu.rf_ram.memory[545][1] ;
 wire \mod.u_cpu.rf_ram.memory[546][0] ;
 wire \mod.u_cpu.rf_ram.memory[546][1] ;
 wire \mod.u_cpu.rf_ram.memory[547][0] ;
 wire \mod.u_cpu.rf_ram.memory[547][1] ;
 wire \mod.u_cpu.rf_ram.memory[548][0] ;
 wire \mod.u_cpu.rf_ram.memory[548][1] ;
 wire \mod.u_cpu.rf_ram.memory[549][0] ;
 wire \mod.u_cpu.rf_ram.memory[549][1] ;
 wire \mod.u_cpu.rf_ram.memory[54][0] ;
 wire \mod.u_cpu.rf_ram.memory[54][1] ;
 wire \mod.u_cpu.rf_ram.memory[550][0] ;
 wire \mod.u_cpu.rf_ram.memory[550][1] ;
 wire \mod.u_cpu.rf_ram.memory[551][0] ;
 wire \mod.u_cpu.rf_ram.memory[551][1] ;
 wire \mod.u_cpu.rf_ram.memory[552][0] ;
 wire \mod.u_cpu.rf_ram.memory[552][1] ;
 wire \mod.u_cpu.rf_ram.memory[553][0] ;
 wire \mod.u_cpu.rf_ram.memory[553][1] ;
 wire \mod.u_cpu.rf_ram.memory[554][0] ;
 wire \mod.u_cpu.rf_ram.memory[554][1] ;
 wire \mod.u_cpu.rf_ram.memory[555][0] ;
 wire \mod.u_cpu.rf_ram.memory[555][1] ;
 wire \mod.u_cpu.rf_ram.memory[556][0] ;
 wire \mod.u_cpu.rf_ram.memory[556][1] ;
 wire \mod.u_cpu.rf_ram.memory[557][0] ;
 wire \mod.u_cpu.rf_ram.memory[557][1] ;
 wire \mod.u_cpu.rf_ram.memory[558][0] ;
 wire \mod.u_cpu.rf_ram.memory[558][1] ;
 wire \mod.u_cpu.rf_ram.memory[559][0] ;
 wire \mod.u_cpu.rf_ram.memory[559][1] ;
 wire \mod.u_cpu.rf_ram.memory[55][0] ;
 wire \mod.u_cpu.rf_ram.memory[55][1] ;
 wire \mod.u_cpu.rf_ram.memory[560][0] ;
 wire \mod.u_cpu.rf_ram.memory[560][1] ;
 wire \mod.u_cpu.rf_ram.memory[561][0] ;
 wire \mod.u_cpu.rf_ram.memory[561][1] ;
 wire \mod.u_cpu.rf_ram.memory[562][0] ;
 wire \mod.u_cpu.rf_ram.memory[562][1] ;
 wire \mod.u_cpu.rf_ram.memory[563][0] ;
 wire \mod.u_cpu.rf_ram.memory[563][1] ;
 wire \mod.u_cpu.rf_ram.memory[564][0] ;
 wire \mod.u_cpu.rf_ram.memory[564][1] ;
 wire \mod.u_cpu.rf_ram.memory[565][0] ;
 wire \mod.u_cpu.rf_ram.memory[565][1] ;
 wire \mod.u_cpu.rf_ram.memory[566][0] ;
 wire \mod.u_cpu.rf_ram.memory[566][1] ;
 wire \mod.u_cpu.rf_ram.memory[567][0] ;
 wire \mod.u_cpu.rf_ram.memory[567][1] ;
 wire \mod.u_cpu.rf_ram.memory[568][0] ;
 wire \mod.u_cpu.rf_ram.memory[568][1] ;
 wire \mod.u_cpu.rf_ram.memory[569][0] ;
 wire \mod.u_cpu.rf_ram.memory[569][1] ;
 wire \mod.u_cpu.rf_ram.memory[56][0] ;
 wire \mod.u_cpu.rf_ram.memory[56][1] ;
 wire \mod.u_cpu.rf_ram.memory[570][0] ;
 wire \mod.u_cpu.rf_ram.memory[570][1] ;
 wire \mod.u_cpu.rf_ram.memory[571][0] ;
 wire \mod.u_cpu.rf_ram.memory[571][1] ;
 wire \mod.u_cpu.rf_ram.memory[572][0] ;
 wire \mod.u_cpu.rf_ram.memory[572][1] ;
 wire \mod.u_cpu.rf_ram.memory[573][0] ;
 wire \mod.u_cpu.rf_ram.memory[573][1] ;
 wire \mod.u_cpu.rf_ram.memory[574][0] ;
 wire \mod.u_cpu.rf_ram.memory[574][1] ;
 wire \mod.u_cpu.rf_ram.memory[575][0] ;
 wire \mod.u_cpu.rf_ram.memory[575][1] ;
 wire \mod.u_cpu.rf_ram.memory[57][0] ;
 wire \mod.u_cpu.rf_ram.memory[57][1] ;
 wire \mod.u_cpu.rf_ram.memory[58][0] ;
 wire \mod.u_cpu.rf_ram.memory[58][1] ;
 wire \mod.u_cpu.rf_ram.memory[59][0] ;
 wire \mod.u_cpu.rf_ram.memory[59][1] ;
 wire \mod.u_cpu.rf_ram.memory[5][0] ;
 wire \mod.u_cpu.rf_ram.memory[5][1] ;
 wire \mod.u_cpu.rf_ram.memory[60][0] ;
 wire \mod.u_cpu.rf_ram.memory[60][1] ;
 wire \mod.u_cpu.rf_ram.memory[61][0] ;
 wire \mod.u_cpu.rf_ram.memory[61][1] ;
 wire \mod.u_cpu.rf_ram.memory[62][0] ;
 wire \mod.u_cpu.rf_ram.memory[62][1] ;
 wire \mod.u_cpu.rf_ram.memory[63][0] ;
 wire \mod.u_cpu.rf_ram.memory[63][1] ;
 wire \mod.u_cpu.rf_ram.memory[64][0] ;
 wire \mod.u_cpu.rf_ram.memory[64][1] ;
 wire \mod.u_cpu.rf_ram.memory[65][0] ;
 wire \mod.u_cpu.rf_ram.memory[65][1] ;
 wire \mod.u_cpu.rf_ram.memory[66][0] ;
 wire \mod.u_cpu.rf_ram.memory[66][1] ;
 wire \mod.u_cpu.rf_ram.memory[67][0] ;
 wire \mod.u_cpu.rf_ram.memory[67][1] ;
 wire \mod.u_cpu.rf_ram.memory[68][0] ;
 wire \mod.u_cpu.rf_ram.memory[68][1] ;
 wire \mod.u_cpu.rf_ram.memory[69][0] ;
 wire \mod.u_cpu.rf_ram.memory[69][1] ;
 wire \mod.u_cpu.rf_ram.memory[6][0] ;
 wire \mod.u_cpu.rf_ram.memory[6][1] ;
 wire \mod.u_cpu.rf_ram.memory[70][0] ;
 wire \mod.u_cpu.rf_ram.memory[70][1] ;
 wire \mod.u_cpu.rf_ram.memory[71][0] ;
 wire \mod.u_cpu.rf_ram.memory[71][1] ;
 wire \mod.u_cpu.rf_ram.memory[72][0] ;
 wire \mod.u_cpu.rf_ram.memory[72][1] ;
 wire \mod.u_cpu.rf_ram.memory[73][0] ;
 wire \mod.u_cpu.rf_ram.memory[73][1] ;
 wire \mod.u_cpu.rf_ram.memory[74][0] ;
 wire \mod.u_cpu.rf_ram.memory[74][1] ;
 wire \mod.u_cpu.rf_ram.memory[75][0] ;
 wire \mod.u_cpu.rf_ram.memory[75][1] ;
 wire \mod.u_cpu.rf_ram.memory[76][0] ;
 wire \mod.u_cpu.rf_ram.memory[76][1] ;
 wire \mod.u_cpu.rf_ram.memory[77][0] ;
 wire \mod.u_cpu.rf_ram.memory[77][1] ;
 wire \mod.u_cpu.rf_ram.memory[78][0] ;
 wire \mod.u_cpu.rf_ram.memory[78][1] ;
 wire \mod.u_cpu.rf_ram.memory[79][0] ;
 wire \mod.u_cpu.rf_ram.memory[79][1] ;
 wire \mod.u_cpu.rf_ram.memory[7][0] ;
 wire \mod.u_cpu.rf_ram.memory[7][1] ;
 wire \mod.u_cpu.rf_ram.memory[80][0] ;
 wire \mod.u_cpu.rf_ram.memory[80][1] ;
 wire \mod.u_cpu.rf_ram.memory[81][0] ;
 wire \mod.u_cpu.rf_ram.memory[81][1] ;
 wire \mod.u_cpu.rf_ram.memory[82][0] ;
 wire \mod.u_cpu.rf_ram.memory[82][1] ;
 wire \mod.u_cpu.rf_ram.memory[83][0] ;
 wire \mod.u_cpu.rf_ram.memory[83][1] ;
 wire \mod.u_cpu.rf_ram.memory[84][0] ;
 wire \mod.u_cpu.rf_ram.memory[84][1] ;
 wire \mod.u_cpu.rf_ram.memory[85][0] ;
 wire \mod.u_cpu.rf_ram.memory[85][1] ;
 wire \mod.u_cpu.rf_ram.memory[86][0] ;
 wire \mod.u_cpu.rf_ram.memory[86][1] ;
 wire \mod.u_cpu.rf_ram.memory[87][0] ;
 wire \mod.u_cpu.rf_ram.memory[87][1] ;
 wire \mod.u_cpu.rf_ram.memory[88][0] ;
 wire \mod.u_cpu.rf_ram.memory[88][1] ;
 wire \mod.u_cpu.rf_ram.memory[89][0] ;
 wire \mod.u_cpu.rf_ram.memory[89][1] ;
 wire \mod.u_cpu.rf_ram.memory[8][0] ;
 wire \mod.u_cpu.rf_ram.memory[8][1] ;
 wire \mod.u_cpu.rf_ram.memory[90][0] ;
 wire \mod.u_cpu.rf_ram.memory[90][1] ;
 wire \mod.u_cpu.rf_ram.memory[91][0] ;
 wire \mod.u_cpu.rf_ram.memory[91][1] ;
 wire \mod.u_cpu.rf_ram.memory[92][0] ;
 wire \mod.u_cpu.rf_ram.memory[92][1] ;
 wire \mod.u_cpu.rf_ram.memory[93][0] ;
 wire \mod.u_cpu.rf_ram.memory[93][1] ;
 wire \mod.u_cpu.rf_ram.memory[94][0] ;
 wire \mod.u_cpu.rf_ram.memory[94][1] ;
 wire \mod.u_cpu.rf_ram.memory[95][0] ;
 wire \mod.u_cpu.rf_ram.memory[95][1] ;
 wire \mod.u_cpu.rf_ram.memory[96][0] ;
 wire \mod.u_cpu.rf_ram.memory[96][1] ;
 wire \mod.u_cpu.rf_ram.memory[97][0] ;
 wire \mod.u_cpu.rf_ram.memory[97][1] ;
 wire \mod.u_cpu.rf_ram.memory[98][0] ;
 wire \mod.u_cpu.rf_ram.memory[98][1] ;
 wire \mod.u_cpu.rf_ram.memory[99][0] ;
 wire \mod.u_cpu.rf_ram.memory[99][1] ;
 wire \mod.u_cpu.rf_ram.memory[9][0] ;
 wire \mod.u_cpu.rf_ram.memory[9][1] ;
 wire \mod.u_cpu.rf_ram.rdata[0] ;
 wire \mod.u_cpu.rf_ram.rdata[1] ;
 wire \mod.u_cpu.rf_ram.regzero ;
 wire \mod.u_cpu.rf_ram_if.rdata0[1] ;
 wire \mod.u_cpu.rf_ram_if.rdata1 ;
 wire \mod.u_cpu.rf_ram_if.rgnt ;
 wire \mod.u_cpu.rf_ram_if.rreq_r ;
 wire \mod.u_cpu.rf_ram_if.rtrig0 ;
 wire \mod.u_cpu.rf_ram_if.rtrig1 ;
 wire \mod.u_cpu.rf_ram_if.wdata0_r ;
 wire \mod.u_cpu.rf_ram_if.wdata1_r[0] ;
 wire \mod.u_cpu.rf_ram_if.wdata1_r[1] ;
 wire \mod.u_cpu.rf_ram_if.wen0_r ;
 wire \mod.u_cpu.rf_ram_if.wen1_r ;
 wire \mod.u_scanchain_local.module_data_in[34] ;
 wire \mod.u_scanchain_local.module_data_in[35] ;
 wire \mod.u_scanchain_local.module_data_in[36] ;
 wire \mod.u_scanchain_local.module_data_in[37] ;
 wire \mod.u_scanchain_local.module_data_in[38] ;
 wire \mod.u_scanchain_local.module_data_in[39] ;
 wire \mod.u_scanchain_local.module_data_in[40] ;
 wire \mod.u_scanchain_local.module_data_in[41] ;
 wire \mod.u_scanchain_local.module_data_in[42] ;
 wire \mod.u_scanchain_local.module_data_in[43] ;
 wire \mod.u_scanchain_local.module_data_in[44] ;
 wire \mod.u_scanchain_local.module_data_in[45] ;
 wire \mod.u_scanchain_local.module_data_in[46] ;
 wire \mod.u_scanchain_local.module_data_in[47] ;
 wire \mod.u_scanchain_local.module_data_in[48] ;
 wire \mod.u_scanchain_local.module_data_in[49] ;
 wire \mod.u_scanchain_local.module_data_in[50] ;
 wire \mod.u_scanchain_local.module_data_in[51] ;
 wire \mod.u_scanchain_local.module_data_in[52] ;
 wire \mod.u_scanchain_local.module_data_in[53] ;
 wire \mod.u_scanchain_local.module_data_in[54] ;
 wire \mod.u_scanchain_local.module_data_in[55] ;
 wire \mod.u_scanchain_local.module_data_in[56] ;
 wire \mod.u_scanchain_local.module_data_in[57] ;
 wire \mod.u_scanchain_local.module_data_in[58] ;
 wire \mod.u_scanchain_local.module_data_in[59] ;
 wire \mod.u_scanchain_local.module_data_in[60] ;
 wire \mod.u_scanchain_local.module_data_in[61] ;
 wire \mod.u_scanchain_local.module_data_in[62] ;
 wire \mod.u_scanchain_local.module_data_in[63] ;
 wire \mod.u_scanchain_local.module_data_in[64] ;
 wire \mod.u_scanchain_local.module_data_in[65] ;
 wire \mod.u_scanchain_local.module_data_in[66] ;
 wire \mod.u_scanchain_local.module_data_in[67] ;
 wire \mod.u_scanchain_local.module_data_in[68] ;
 wire \mod.u_scanchain_local.module_data_in[69] ;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net152;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net153;
 wire net181;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;

 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07109_ (.I(\mod.u_cpu.rf_ram_if.rtrig0 ),
    .Z(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07110_ (.A1(_01418_),
    .A2(\mod.u_cpu.cpu.csr_imm ),
    .ZN(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07111_ (.A1(\mod.u_cpu.cpu.decode.co_mem_word ),
    .A2(\mod.u_cpu.cpu.bne_or_bge ),
    .A3(\mod.u_cpu.cpu.csr_d_sel ),
    .ZN(_01420_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07112_ (.I(\mod.u_cpu.cpu.decode.opcode[2] ),
    .Z(_01421_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07113_ (.I(\mod.u_cpu.cpu.branch_op ),
    .Z(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07114_ (.A1(_01421_),
    .A2(_01422_),
    .Z(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07115_ (.I(_01423_),
    .Z(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07116_ (.A1(\mod.u_cpu.cpu.decode.op21 ),
    .A2(_01420_),
    .A3(_01424_),
    .ZN(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07117_ (.I(\mod.u_cpu.cpu.decode.op26 ),
    .ZN(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07118_ (.A1(\mod.u_cpu.cpu.decode.op21 ),
    .A2(_01426_),
    .ZN(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07119_ (.I(\mod.u_cpu.cpu.decode.co_mem_word ),
    .Z(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07120_ (.I(\mod.u_cpu.cpu.bne_or_bge ),
    .Z(_01429_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07121_ (.I(\mod.u_cpu.cpu.csr_d_sel ),
    .Z(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _07122_ (.A1(_01428_),
    .A2(_01429_),
    .A3(_01430_),
    .Z(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07123_ (.A1(\mod.u_cpu.cpu.decode.co_ebreak ),
    .A2(_01427_),
    .B(_01424_),
    .C(_01431_),
    .ZN(_01432_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07124_ (.I(\mod.u_cpu.cpu.state.genblk1.misalign_trap_sync_r ),
    .Z(_01433_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07125_ (.I(\mod.u_cpu.cpu.genblk3.csr.o_new_irq ),
    .Z(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07126_ (.I(\mod.u_cpu.cpu.decode.op21 ),
    .ZN(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07127_ (.A1(_01435_),
    .A2(_01420_),
    .A3(_01423_),
    .Z(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07128_ (.A1(_01433_),
    .A2(_01434_),
    .A3(_01436_),
    .ZN(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07129_ (.A1(_01425_),
    .A2(_01432_),
    .A3(_01437_),
    .Z(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07130_ (.I(\mod.u_cpu.rf_ram_if.rtrig0 ),
    .Z(_01439_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07131_ (.I(_01437_),
    .Z(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07132_ (.A1(_01439_),
    .A2(_01440_),
    .ZN(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07133_ (.A1(_01427_),
    .A2(_01432_),
    .ZN(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07134_ (.A1(\mod.u_cpu.cpu.immdec.imm24_20[0] ),
    .A2(_01438_),
    .B(_01441_),
    .C(_01442_),
    .ZN(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07135_ (.A1(_01419_),
    .A2(_01443_),
    .ZN(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07136_ (.I(_01444_),
    .Z(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07137_ (.I(_01445_),
    .Z(_01446_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07138_ (.I(_01446_),
    .Z(_01447_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07139_ (.I(_01439_),
    .Z(_01448_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07140_ (.I(_01448_),
    .Z(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07141_ (.A1(_01449_),
    .A2(\mod.u_cpu.cpu.immdec.imm19_12_20[5] ),
    .ZN(_01450_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07142_ (.A1(_01432_),
    .A2(_01440_),
    .Z(_01451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07143_ (.A1(_01431_),
    .A2(_01423_),
    .ZN(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07144_ (.I(\mod.u_cpu.cpu.decode.co_ebreak ),
    .Z(_01453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07145_ (.A1(\mod.u_cpu.cpu.decode.op26 ),
    .A2(_01453_),
    .ZN(_01454_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07146_ (.A1(_01452_),
    .A2(_01454_),
    .B(_01448_),
    .C(_01425_),
    .ZN(_01455_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07147_ (.A1(\mod.u_cpu.cpu.immdec.imm24_20[1] ),
    .A2(_01451_),
    .B(_01455_),
    .ZN(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07148_ (.A1(_01450_),
    .A2(_01456_),
    .ZN(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07149_ (.I(_01457_),
    .Z(_01458_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07150_ (.I(_01458_),
    .Z(_01459_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07151_ (.I(_01439_),
    .ZN(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07152_ (.I(_01460_),
    .Z(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07153_ (.I(_01461_),
    .Z(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07154_ (.I(_01462_),
    .Z(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07155_ (.I(_01463_),
    .Z(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07156_ (.I(_01438_),
    .Z(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07157_ (.A1(_01464_),
    .A2(_01465_),
    .ZN(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07158_ (.A1(_01449_),
    .A2(_01465_),
    .Z(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07159_ (.A1(_01463_),
    .A2(\mod.u_cpu.cpu.immdec.imm19_12_20[8] ),
    .B1(_01467_),
    .B2(\mod.u_cpu.cpu.immdec.imm24_20[4] ),
    .ZN(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07160_ (.I(_01468_),
    .Z(_01469_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07161_ (.A1(_01463_),
    .A2(\mod.u_cpu.cpu.immdec.imm19_12_20[7] ),
    .B1(_01467_),
    .B2(\mod.u_cpu.cpu.immdec.imm24_20[3] ),
    .ZN(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07162_ (.I(_01470_),
    .Z(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07163_ (.A1(\mod.u_cpu.cpu.immdec.imm24_20[2] ),
    .A2(_01467_),
    .ZN(_01472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07164_ (.A1(_01462_),
    .A2(\mod.u_cpu.cpu.immdec.imm19_12_20[6] ),
    .ZN(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07165_ (.A1(_01472_),
    .A2(_01473_),
    .Z(_01474_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07166_ (.I(_01474_),
    .Z(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07167_ (.A1(_01469_),
    .A2(_01471_),
    .A3(_01475_),
    .ZN(_01476_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _07168_ (.A1(_01447_),
    .A2(_01459_),
    .A3(_01466_),
    .A4(_01476_),
    .ZN(_01477_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07169_ (.I(_01477_),
    .Z(_00007_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07170_ (.I(_01449_),
    .Z(_01478_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07171_ (.I(\mod.u_cpu.cpu.immdec.imm19_12_20[7] ),
    .ZN(_01479_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07172_ (.A1(\mod.u_cpu.cpu.immdec.imm24_20[3] ),
    .A2(_01467_),
    .ZN(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07173_ (.A1(_01478_),
    .A2(_01479_),
    .B(_01480_),
    .ZN(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07174_ (.A1(_01472_),
    .A2(_01473_),
    .ZN(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07175_ (.I(_01482_),
    .Z(_01483_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07176_ (.A1(_01450_),
    .A2(_01456_),
    .Z(_01484_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07177_ (.I(_01484_),
    .Z(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07178_ (.I(_01485_),
    .Z(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07179_ (.A1(_01419_),
    .A2(_01443_),
    .Z(_01487_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07180_ (.I(_01487_),
    .Z(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07181_ (.I(_01488_),
    .Z(_01489_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07182_ (.I(\mod.u_cpu.raddr[2] ),
    .Z(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07183_ (.I(_01490_),
    .Z(_01491_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07184_ (.I(_01491_),
    .Z(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07185_ (.I(_01492_),
    .Z(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07186_ (.I(\mod.u_cpu.raddr[0] ),
    .Z(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07187_ (.I(_01494_),
    .Z(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07188_ (.I(_01495_),
    .Z(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07189_ (.I(\mod.u_cpu.raddr[1] ),
    .Z(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07190_ (.I(_01497_),
    .Z(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07191_ (.I(_01498_),
    .Z(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07192_ (.I(_01499_),
    .Z(_01500_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07193_ (.I(_01500_),
    .Z(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07194_ (.I0(\mod.u_cpu.rf_ram.memory[448][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[449][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[450][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[451][0] ),
    .S0(_01496_),
    .S1(_01501_),
    .Z(_01502_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07195_ (.I(_01498_),
    .Z(_01503_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07196_ (.I(_01503_),
    .Z(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07197_ (.I(_01504_),
    .Z(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07198_ (.I(\mod.u_cpu.raddr[0] ),
    .Z(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07199_ (.I(_01506_),
    .Z(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07200_ (.I(_01507_),
    .Z(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07201_ (.I(_01506_),
    .Z(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07202_ (.I(_01509_),
    .Z(_01510_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07203_ (.I(_01510_),
    .Z(_01511_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07204_ (.I(\mod.u_cpu.rf_ram.memory[453][0] ),
    .ZN(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07205_ (.A1(_01511_),
    .A2(_01512_),
    .ZN(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07206_ (.A1(_01508_),
    .A2(\mod.u_cpu.rf_ram.memory[452][0] ),
    .B(_01513_),
    .ZN(_01514_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07207_ (.I(\mod.u_cpu.raddr[0] ),
    .Z(_01515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07208_ (.I(_01515_),
    .Z(_01516_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07209_ (.I(_01516_),
    .Z(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07210_ (.I(_01515_),
    .Z(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07211_ (.I(_01518_),
    .Z(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07212_ (.I(_01519_),
    .Z(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07213_ (.I(\mod.u_cpu.rf_ram.memory[455][0] ),
    .ZN(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07214_ (.A1(_01520_),
    .A2(_01521_),
    .ZN(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07215_ (.I(_01497_),
    .Z(_01523_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07216_ (.I(_01523_),
    .Z(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07217_ (.I(_01524_),
    .Z(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07218_ (.A1(_01517_),
    .A2(\mod.u_cpu.rf_ram.memory[454][0] ),
    .B(_01522_),
    .C(_01525_),
    .ZN(_01526_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07219_ (.I(_01490_),
    .Z(_01527_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07220_ (.I(_01527_),
    .Z(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07221_ (.I(_01528_),
    .Z(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07222_ (.A1(_01505_),
    .A2(_01514_),
    .B(_01526_),
    .C(_01529_),
    .ZN(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07223_ (.I(\mod.u_cpu.raddr[3] ),
    .ZN(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07224_ (.I(_01531_),
    .Z(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07225_ (.I(_01532_),
    .Z(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07226_ (.I(_01533_),
    .Z(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07227_ (.A1(_01493_),
    .A2(_01502_),
    .B(_01530_),
    .C(_01534_),
    .ZN(_01535_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07228_ (.I(_01492_),
    .Z(_01536_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07229_ (.I(_01515_),
    .Z(_01537_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07230_ (.I(_01537_),
    .Z(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07231_ (.I(_01538_),
    .Z(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07232_ (.I(_01539_),
    .Z(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07233_ (.I0(\mod.u_cpu.rf_ram.memory[456][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[457][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[458][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[459][0] ),
    .S0(_01540_),
    .S1(_01501_),
    .Z(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07234_ (.I(\mod.u_cpu.rf_ram.memory[461][0] ),
    .ZN(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07235_ (.A1(_01511_),
    .A2(_01542_),
    .ZN(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07236_ (.A1(_01508_),
    .A2(\mod.u_cpu.rf_ram.memory[460][0] ),
    .B(_01543_),
    .ZN(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07237_ (.I(_01516_),
    .Z(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07238_ (.I(\mod.u_cpu.rf_ram.memory[463][0] ),
    .ZN(_01546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07239_ (.A1(_01520_),
    .A2(_01546_),
    .ZN(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07240_ (.A1(_01545_),
    .A2(\mod.u_cpu.rf_ram.memory[462][0] ),
    .B(_01547_),
    .C(_01525_),
    .ZN(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07241_ (.A1(_01505_),
    .A2(_01544_),
    .B(_01548_),
    .C(_01529_),
    .ZN(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07242_ (.I(\mod.u_cpu.raddr[3] ),
    .Z(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07243_ (.I(_01550_),
    .Z(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07244_ (.I(_01551_),
    .Z(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07245_ (.A1(_01536_),
    .A2(_01541_),
    .B(_01549_),
    .C(_01552_),
    .ZN(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07246_ (.A1(_01489_),
    .A2(_01535_),
    .A3(_01553_),
    .ZN(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07247_ (.I0(\mod.u_cpu.rf_ram.memory[472][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[473][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[474][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[475][0] ),
    .S0(_01540_),
    .S1(_01501_),
    .Z(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07248_ (.I(_01539_),
    .Z(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07249_ (.I(\mod.u_cpu.rf_ram.memory[477][0] ),
    .ZN(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07250_ (.A1(_01511_),
    .A2(_01557_),
    .ZN(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07251_ (.A1(_01556_),
    .A2(\mod.u_cpu.rf_ram.memory[476][0] ),
    .B(_01558_),
    .ZN(_01559_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07252_ (.I(\mod.u_cpu.raddr[0] ),
    .Z(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07253_ (.I(_01560_),
    .Z(_01561_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07254_ (.I(\mod.u_cpu.rf_ram.memory[479][0] ),
    .ZN(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07255_ (.A1(_01561_),
    .A2(_01562_),
    .ZN(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07256_ (.A1(_01545_),
    .A2(\mod.u_cpu.rf_ram.memory[478][0] ),
    .B(_01563_),
    .C(_01525_),
    .ZN(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07257_ (.A1(_01505_),
    .A2(_01559_),
    .B(_01564_),
    .C(_01529_),
    .ZN(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07258_ (.A1(_01536_),
    .A2(_01555_),
    .B(_01565_),
    .C(_01552_),
    .ZN(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07259_ (.I(_01495_),
    .Z(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07260_ (.I(_01497_),
    .Z(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07261_ (.I(_01568_),
    .Z(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07262_ (.I(_01569_),
    .Z(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07263_ (.I0(\mod.u_cpu.rf_ram.memory[464][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[465][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[466][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[467][0] ),
    .S0(_01567_),
    .S1(_01570_),
    .Z(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07264_ (.I(_01504_),
    .Z(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07265_ (.I(_01510_),
    .Z(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07266_ (.I(\mod.u_cpu.rf_ram.memory[469][0] ),
    .ZN(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07267_ (.A1(_01573_),
    .A2(_01574_),
    .ZN(_01575_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07268_ (.A1(_01556_),
    .A2(\mod.u_cpu.rf_ram.memory[468][0] ),
    .B(_01575_),
    .ZN(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07269_ (.I(_01516_),
    .Z(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07270_ (.I(_01560_),
    .Z(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07271_ (.I(\mod.u_cpu.rf_ram.memory[471][0] ),
    .ZN(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07272_ (.A1(_01578_),
    .A2(_01579_),
    .ZN(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07273_ (.I(_01523_),
    .Z(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07274_ (.I(_01581_),
    .Z(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07275_ (.A1(_01577_),
    .A2(\mod.u_cpu.rf_ram.memory[470][0] ),
    .B(_01580_),
    .C(_01582_),
    .ZN(_01583_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07276_ (.I(_01528_),
    .Z(_01584_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07277_ (.A1(_01572_),
    .A2(_01576_),
    .B(_01583_),
    .C(_01584_),
    .ZN(_01585_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07278_ (.I(_01532_),
    .Z(_01586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07279_ (.I(_01586_),
    .Z(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07280_ (.A1(_01536_),
    .A2(_01571_),
    .B(_01585_),
    .C(_01587_),
    .ZN(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07281_ (.A1(_01446_),
    .A2(_01566_),
    .A3(_01588_),
    .ZN(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07282_ (.A1(_01486_),
    .A2(_01554_),
    .A3(_01589_),
    .ZN(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07283_ (.I(_01458_),
    .Z(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07284_ (.I(_01445_),
    .Z(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07285_ (.I0(\mod.u_cpu.rf_ram.memory[496][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[497][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[498][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[499][0] ),
    .S0(_01540_),
    .S1(_01570_),
    .Z(_01593_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07286_ (.I(\mod.u_cpu.rf_ram.memory[501][0] ),
    .ZN(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07287_ (.A1(_01573_),
    .A2(_01594_),
    .ZN(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07288_ (.A1(_01556_),
    .A2(\mod.u_cpu.rf_ram.memory[500][0] ),
    .B(_01595_),
    .ZN(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07289_ (.I(\mod.u_cpu.rf_ram.memory[503][0] ),
    .ZN(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07290_ (.A1(_01561_),
    .A2(_01597_),
    .ZN(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07291_ (.A1(_01545_),
    .A2(\mod.u_cpu.rf_ram.memory[502][0] ),
    .B(_01598_),
    .C(_01582_),
    .ZN(_01599_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07292_ (.A1(_01505_),
    .A2(_01596_),
    .B(_01599_),
    .C(_01584_),
    .ZN(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07293_ (.A1(_01536_),
    .A2(_01593_),
    .B(_01600_),
    .C(_01587_),
    .ZN(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07294_ (.I(_01492_),
    .Z(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07295_ (.I(_01495_),
    .Z(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07296_ (.I(_01603_),
    .Z(_01604_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07297_ (.I(_01604_),
    .Z(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07298_ (.I0(\mod.u_cpu.rf_ram.memory[504][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[505][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[506][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[507][0] ),
    .S0(_01605_),
    .S1(_01570_),
    .Z(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07299_ (.I(_01539_),
    .Z(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07300_ (.I(_01510_),
    .Z(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07301_ (.I(\mod.u_cpu.rf_ram.memory[509][0] ),
    .ZN(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07302_ (.A1(_01608_),
    .A2(_01609_),
    .ZN(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07303_ (.A1(_01607_),
    .A2(\mod.u_cpu.rf_ram.memory[508][0] ),
    .B(_01610_),
    .ZN(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07304_ (.I(\mod.u_cpu.rf_ram.memory[511][0] ),
    .ZN(_01612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07305_ (.A1(_01578_),
    .A2(_01612_),
    .ZN(_01613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07306_ (.I(_01523_),
    .Z(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07307_ (.I(_01614_),
    .Z(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07308_ (.A1(_01577_),
    .A2(\mod.u_cpu.rf_ram.memory[510][0] ),
    .B(_01613_),
    .C(_01615_),
    .ZN(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07309_ (.A1(_01572_),
    .A2(_01611_),
    .B(_01616_),
    .C(_01584_),
    .ZN(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07310_ (.I(_01551_),
    .Z(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07311_ (.A1(_01602_),
    .A2(_01606_),
    .B(_01617_),
    .C(_01618_),
    .ZN(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07312_ (.A1(_01592_),
    .A2(_01601_),
    .A3(_01619_),
    .ZN(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07313_ (.I0(\mod.u_cpu.rf_ram.memory[480][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[481][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[482][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[483][0] ),
    .S0(_01605_),
    .S1(_01570_),
    .Z(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07314_ (.I(\mod.u_cpu.rf_ram.memory[485][0] ),
    .ZN(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07315_ (.A1(_01573_),
    .A2(_01622_),
    .ZN(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07316_ (.A1(_01556_),
    .A2(\mod.u_cpu.rf_ram.memory[484][0] ),
    .B(_01623_),
    .ZN(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07317_ (.I(\mod.u_cpu.rf_ram.memory[487][0] ),
    .ZN(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07318_ (.A1(_01578_),
    .A2(_01625_),
    .ZN(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07319_ (.A1(_01577_),
    .A2(\mod.u_cpu.rf_ram.memory[486][0] ),
    .B(_01626_),
    .C(_01582_),
    .ZN(_01627_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07320_ (.A1(_01572_),
    .A2(_01624_),
    .B(_01627_),
    .C(_01584_),
    .ZN(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07321_ (.A1(_01602_),
    .A2(_01621_),
    .B(_01628_),
    .C(_01587_),
    .ZN(_01629_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07322_ (.I(_01490_),
    .Z(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07323_ (.I(_01630_),
    .Z(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07324_ (.I(_01631_),
    .Z(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07325_ (.I(_01494_),
    .Z(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07326_ (.I(_01633_),
    .Z(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07327_ (.I(_01634_),
    .Z(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07328_ (.I(_01635_),
    .Z(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07329_ (.I(_01568_),
    .Z(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07330_ (.I(_01637_),
    .Z(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07331_ (.I0(\mod.u_cpu.rf_ram.memory[488][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[489][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[490][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[491][0] ),
    .S0(_01636_),
    .S1(_01638_),
    .Z(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07332_ (.I(\mod.u_cpu.rf_ram.memory[493][0] ),
    .ZN(_01640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07333_ (.A1(_01608_),
    .A2(_01640_),
    .ZN(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07334_ (.A1(_01607_),
    .A2(\mod.u_cpu.rf_ram.memory[492][0] ),
    .B(_01641_),
    .ZN(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07335_ (.I(_01604_),
    .Z(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07336_ (.I(_01494_),
    .Z(_01644_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07337_ (.I(_01644_),
    .Z(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07338_ (.I(_01645_),
    .Z(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07339_ (.I(_01646_),
    .Z(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07340_ (.I(\mod.u_cpu.rf_ram.memory[495][0] ),
    .ZN(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07341_ (.A1(_01647_),
    .A2(_01648_),
    .ZN(_01649_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07342_ (.A1(_01643_),
    .A2(\mod.u_cpu.rf_ram.memory[494][0] ),
    .B(_01649_),
    .C(_01615_),
    .ZN(_01650_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07343_ (.I(_01528_),
    .Z(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07344_ (.A1(_01572_),
    .A2(_01642_),
    .B(_01650_),
    .C(_01651_),
    .ZN(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07345_ (.A1(_01632_),
    .A2(_01639_),
    .B(_01652_),
    .C(_01618_),
    .ZN(_01653_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07346_ (.A1(_01489_),
    .A2(_01629_),
    .A3(_01653_),
    .ZN(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07347_ (.A1(_01591_),
    .A2(_01620_),
    .A3(_01654_),
    .ZN(_01655_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07348_ (.A1(_01483_),
    .A2(_01590_),
    .A3(_01655_),
    .ZN(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07349_ (.I(_01532_),
    .Z(_01657_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07350_ (.I(_01657_),
    .Z(_01658_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07351_ (.I(\mod.u_cpu.raddr[2] ),
    .ZN(_01659_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07352_ (.I(_01659_),
    .Z(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07353_ (.I(_01660_),
    .Z(_01661_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07354_ (.I(_01661_),
    .Z(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07355_ (.I(_01538_),
    .Z(_01663_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07356_ (.I(_01663_),
    .Z(_01664_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07357_ (.I(_01499_),
    .Z(_01665_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07358_ (.I(_01665_),
    .Z(_01666_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07359_ (.I0(\mod.u_cpu.rf_ram.memory[384][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[385][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[386][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[387][0] ),
    .S0(_01664_),
    .S1(_01666_),
    .Z(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07360_ (.A1(_01662_),
    .A2(_01667_),
    .ZN(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07361_ (.I(_01491_),
    .Z(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07362_ (.I(_01669_),
    .Z(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07363_ (.I(_01537_),
    .Z(_01671_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07364_ (.I(_01671_),
    .Z(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07365_ (.I(_01672_),
    .Z(_01673_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07366_ (.I0(\mod.u_cpu.rf_ram.memory[388][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[389][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[390][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[391][0] ),
    .S0(_01673_),
    .S1(_01666_),
    .Z(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07367_ (.A1(_01670_),
    .A2(_01674_),
    .ZN(_01675_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07368_ (.A1(_01658_),
    .A2(_01668_),
    .A3(_01675_),
    .ZN(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07369_ (.I(_01550_),
    .Z(_01677_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07370_ (.I(_01677_),
    .Z(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07371_ (.I(_01660_),
    .Z(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07372_ (.I(_01679_),
    .Z(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07373_ (.I(_01509_),
    .Z(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07374_ (.I(_01681_),
    .Z(_01682_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07375_ (.I(_01665_),
    .Z(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07376_ (.I0(\mod.u_cpu.rf_ram.memory[392][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[393][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[394][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[395][0] ),
    .S0(_01682_),
    .S1(_01683_),
    .Z(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07377_ (.A1(_01680_),
    .A2(_01684_),
    .ZN(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07378_ (.I(_01527_),
    .Z(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07379_ (.I(_01686_),
    .Z(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07380_ (.I(_01687_),
    .Z(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07381_ (.I(_01633_),
    .Z(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07382_ (.I0(\mod.u_cpu.rf_ram.memory[396][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[397][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[398][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[399][0] ),
    .S0(_01689_),
    .S1(_01683_),
    .Z(_01690_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07383_ (.A1(_01688_),
    .A2(_01690_),
    .ZN(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07384_ (.A1(_01678_),
    .A2(_01685_),
    .A3(_01691_),
    .ZN(_01692_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07385_ (.I(_01445_),
    .Z(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07386_ (.A1(_01676_),
    .A2(_01692_),
    .B(_01693_),
    .ZN(_01694_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07387_ (.I(_01491_),
    .Z(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07388_ (.I(_01695_),
    .Z(_01696_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07389_ (.I(_01633_),
    .Z(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07390_ (.I(_01500_),
    .Z(_01698_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07391_ (.I0(\mod.u_cpu.rf_ram.memory[408][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[409][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[410][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[411][0] ),
    .S0(_01697_),
    .S1(_01698_),
    .Z(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07392_ (.I(_01497_),
    .Z(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07393_ (.I(_01700_),
    .Z(_01701_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07394_ (.I(_01701_),
    .Z(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07395_ (.I(_01702_),
    .Z(_01703_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07396_ (.I(_01538_),
    .Z(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07397_ (.I(_01704_),
    .Z(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07398_ (.I(\mod.u_cpu.rf_ram.memory[413][0] ),
    .ZN(_01706_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07399_ (.A1(_01567_),
    .A2(_01706_),
    .ZN(_01707_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07400_ (.A1(_01705_),
    .A2(\mod.u_cpu.rf_ram.memory[412][0] ),
    .B(_01707_),
    .ZN(_01708_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07401_ (.I(_01516_),
    .Z(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07402_ (.I(_01509_),
    .Z(_01710_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07403_ (.I(_01710_),
    .Z(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07404_ (.I(\mod.u_cpu.rf_ram.memory[415][0] ),
    .ZN(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07405_ (.A1(_01711_),
    .A2(_01712_),
    .ZN(_01713_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07406_ (.I(_01524_),
    .Z(_01714_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07407_ (.A1(_01709_),
    .A2(\mod.u_cpu.rf_ram.memory[414][0] ),
    .B(_01713_),
    .C(_01714_),
    .ZN(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07408_ (.I(_01527_),
    .Z(_01716_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07409_ (.I(_01716_),
    .Z(_01717_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07410_ (.A1(_01703_),
    .A2(_01708_),
    .B(_01715_),
    .C(_01717_),
    .ZN(_01718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07411_ (.I(_01550_),
    .Z(_01719_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07412_ (.I(_01719_),
    .Z(_01720_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07413_ (.A1(_01696_),
    .A2(_01699_),
    .B(_01718_),
    .C(_01720_),
    .ZN(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07414_ (.I(_01633_),
    .Z(_01722_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07415_ (.I(_01500_),
    .Z(_01723_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07416_ (.I0(\mod.u_cpu.rf_ram.memory[400][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[401][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[402][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[403][0] ),
    .S0(_01722_),
    .S1(_01723_),
    .Z(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07417_ (.I(\mod.u_cpu.rf_ram.memory[405][0] ),
    .ZN(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07418_ (.A1(_01605_),
    .A2(_01725_),
    .ZN(_01726_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07419_ (.A1(_01705_),
    .A2(\mod.u_cpu.rf_ram.memory[404][0] ),
    .B(_01726_),
    .ZN(_01727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07420_ (.I(_01604_),
    .Z(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07421_ (.I(_01519_),
    .Z(_01729_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07422_ (.I(\mod.u_cpu.rf_ram.memory[407][0] ),
    .ZN(_01730_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07423_ (.A1(_01729_),
    .A2(_01730_),
    .ZN(_01731_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07424_ (.I(_01614_),
    .Z(_01732_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07425_ (.A1(_01728_),
    .A2(\mod.u_cpu.rf_ram.memory[406][0] ),
    .B(_01731_),
    .C(_01732_),
    .ZN(_01733_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07426_ (.A1(_01703_),
    .A2(_01727_),
    .B(_01733_),
    .C(_01529_),
    .ZN(_01734_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07427_ (.A1(_01493_),
    .A2(_01724_),
    .B(_01734_),
    .C(_01534_),
    .ZN(_01735_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07428_ (.A1(_01446_),
    .A2(_01721_),
    .A3(_01735_),
    .ZN(_01736_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07429_ (.A1(_01486_),
    .A2(_01736_),
    .ZN(_01737_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07430_ (.I(_01474_),
    .Z(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07431_ (.I(_01458_),
    .Z(_01739_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07432_ (.I(_01488_),
    .Z(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07433_ (.I(_01630_),
    .Z(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07434_ (.I(_01741_),
    .Z(_01742_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07435_ (.I(_01560_),
    .Z(_01743_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07436_ (.I(_01743_),
    .Z(_01744_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07437_ (.I(_01744_),
    .Z(_01745_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07438_ (.I(_01568_),
    .Z(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07439_ (.I(_01746_),
    .Z(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07440_ (.I0(\mod.u_cpu.rf_ram.memory[416][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[417][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[418][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[419][0] ),
    .S0(_01745_),
    .S1(_01747_),
    .Z(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07441_ (.I(_01498_),
    .Z(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07442_ (.I(_01749_),
    .Z(_01750_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07443_ (.I(_01750_),
    .Z(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07444_ (.I(_01645_),
    .Z(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07445_ (.I(_01752_),
    .Z(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07446_ (.I(\mod.u_cpu.rf_ram.memory[421][0] ),
    .ZN(_01754_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07447_ (.A1(_01753_),
    .A2(_01754_),
    .ZN(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07448_ (.A1(_01728_),
    .A2(\mod.u_cpu.rf_ram.memory[420][0] ),
    .B(_01755_),
    .ZN(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07449_ (.I(_01515_),
    .Z(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07450_ (.I(_01757_),
    .Z(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07451_ (.I(_01758_),
    .Z(_01759_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07452_ (.I(\mod.u_cpu.rf_ram.memory[423][0] ),
    .ZN(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07453_ (.A1(_01759_),
    .A2(_01760_),
    .ZN(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07454_ (.I(_01700_),
    .Z(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07455_ (.I(_01762_),
    .Z(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07456_ (.A1(_01689_),
    .A2(\mod.u_cpu.rf_ram.memory[422][0] ),
    .B(_01761_),
    .C(_01763_),
    .ZN(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07457_ (.I(_01527_),
    .Z(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07458_ (.I(_01765_),
    .Z(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07459_ (.A1(_01751_),
    .A2(_01756_),
    .B(_01764_),
    .C(_01766_),
    .ZN(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07460_ (.I(_01586_),
    .Z(_01768_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07461_ (.A1(_01742_),
    .A2(_01748_),
    .B(_01767_),
    .C(_01768_),
    .ZN(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07462_ (.I(_01741_),
    .Z(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07463_ (.I(_01569_),
    .Z(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07464_ (.I0(\mod.u_cpu.rf_ram.memory[424][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[425][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[426][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[427][0] ),
    .S0(_01753_),
    .S1(_01771_),
    .Z(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07465_ (.I(_01750_),
    .Z(_01773_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07466_ (.I(_01744_),
    .Z(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07467_ (.I(\mod.u_cpu.rf_ram.memory[429][0] ),
    .ZN(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07468_ (.A1(_01774_),
    .A2(_01775_),
    .ZN(_01776_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07469_ (.A1(_01728_),
    .A2(\mod.u_cpu.rf_ram.memory[428][0] ),
    .B(_01776_),
    .ZN(_01777_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07470_ (.I(_01757_),
    .Z(_01778_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07471_ (.I(_01778_),
    .Z(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07472_ (.I(\mod.u_cpu.rf_ram.memory[431][0] ),
    .ZN(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07473_ (.A1(_01779_),
    .A2(_01780_),
    .ZN(_01781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07474_ (.I(_01700_),
    .Z(_01782_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07475_ (.I(_01782_),
    .Z(_01783_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07476_ (.A1(_01689_),
    .A2(\mod.u_cpu.rf_ram.memory[430][0] ),
    .B(_01781_),
    .C(_01783_),
    .ZN(_01784_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07477_ (.I(_01765_),
    .Z(_01785_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07478_ (.A1(_01773_),
    .A2(_01777_),
    .B(_01784_),
    .C(_01785_),
    .ZN(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07479_ (.I(\mod.u_cpu.raddr[3] ),
    .Z(_01787_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07480_ (.I(_01787_),
    .Z(_01788_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07481_ (.A1(_01770_),
    .A2(_01772_),
    .B(_01786_),
    .C(_01788_),
    .ZN(_01789_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07482_ (.A1(_01740_),
    .A2(_01769_),
    .A3(_01789_),
    .ZN(_01790_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07483_ (.I(_01445_),
    .Z(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07484_ (.I0(\mod.u_cpu.rf_ram.memory[432][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[433][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[434][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[435][0] ),
    .S0(_01745_),
    .S1(_01747_),
    .Z(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07485_ (.I(\mod.u_cpu.rf_ram.memory[437][0] ),
    .ZN(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07486_ (.A1(_01774_),
    .A2(_01793_),
    .ZN(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07487_ (.A1(_01728_),
    .A2(\mod.u_cpu.rf_ram.memory[436][0] ),
    .B(_01794_),
    .ZN(_01795_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07488_ (.I(\mod.u_cpu.rf_ram.memory[439][0] ),
    .ZN(_01796_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07489_ (.A1(_01779_),
    .A2(_01796_),
    .ZN(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07490_ (.A1(_01689_),
    .A2(\mod.u_cpu.rf_ram.memory[438][0] ),
    .B(_01797_),
    .C(_01763_),
    .ZN(_01798_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07491_ (.A1(_01773_),
    .A2(_01795_),
    .B(_01798_),
    .C(_01785_),
    .ZN(_01799_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07492_ (.A1(_01770_),
    .A2(_01792_),
    .B(_01799_),
    .C(_01768_),
    .ZN(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07493_ (.I0(\mod.u_cpu.rf_ram.memory[440][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[441][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[442][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[443][0] ),
    .S0(_01753_),
    .S1(_01771_),
    .Z(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07494_ (.I(_01752_),
    .Z(_01802_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07495_ (.I(\mod.u_cpu.rf_ram.memory[445][0] ),
    .ZN(_01803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07496_ (.A1(_01802_),
    .A2(_01803_),
    .ZN(_01804_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07497_ (.A1(_01517_),
    .A2(\mod.u_cpu.rf_ram.memory[444][0] ),
    .B(_01804_),
    .ZN(_01805_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07498_ (.I(_01603_),
    .Z(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07499_ (.I(_01806_),
    .Z(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07500_ (.I(\mod.u_cpu.rf_ram.memory[447][0] ),
    .ZN(_01808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07501_ (.A1(_01779_),
    .A2(_01808_),
    .ZN(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07502_ (.A1(_01807_),
    .A2(\mod.u_cpu.rf_ram.memory[446][0] ),
    .B(_01809_),
    .C(_01783_),
    .ZN(_01810_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07503_ (.A1(_01773_),
    .A2(_01805_),
    .B(_01810_),
    .C(_01785_),
    .ZN(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07504_ (.I(_01787_),
    .Z(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07505_ (.A1(_01770_),
    .A2(_01801_),
    .B(_01811_),
    .C(_01812_),
    .ZN(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07506_ (.A1(_01791_),
    .A2(_01800_),
    .A3(_01813_),
    .ZN(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07507_ (.A1(_01739_),
    .A2(_01790_),
    .A3(_01814_),
    .ZN(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07508_ (.A1(_01694_),
    .A2(_01737_),
    .B(_01738_),
    .C(_01815_),
    .ZN(_01816_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07509_ (.A1(_01656_),
    .A2(_01816_),
    .Z(_01817_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07510_ (.I(_01657_),
    .Z(_01818_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07511_ (.I(_01506_),
    .Z(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07512_ (.I(_01523_),
    .Z(_01820_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07513_ (.I(_01820_),
    .Z(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07514_ (.I0(\mod.u_cpu.rf_ram.memory[332][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[333][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[334][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[335][0] ),
    .S0(_01819_),
    .S1(_01821_),
    .Z(_01822_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07515_ (.I(_01506_),
    .Z(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07516_ (.I0(\mod.u_cpu.rf_ram.memory[348][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[349][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[350][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[351][0] ),
    .S0(_01823_),
    .S1(_01821_),
    .Z(_01824_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07517_ (.I(_01743_),
    .Z(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07518_ (.I(_01825_),
    .Z(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07519_ (.I(_01700_),
    .Z(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07520_ (.I(_01827_),
    .Z(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07521_ (.I0(\mod.u_cpu.rf_ram.memory[328][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[329][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[330][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[331][0] ),
    .S0(_01826_),
    .S1(_01828_),
    .Z(_01829_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07522_ (.I(_01820_),
    .Z(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07523_ (.I0(\mod.u_cpu.rf_ram.memory[344][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[345][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[346][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[347][0] ),
    .S0(_01826_),
    .S1(_01830_),
    .Z(_01831_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07524_ (.I(_01444_),
    .Z(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07525_ (.I(_01679_),
    .Z(_01833_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07526_ (.I0(_01822_),
    .I1(_01824_),
    .I2(_01829_),
    .I3(_01831_),
    .S0(_01832_),
    .S1(_01833_),
    .Z(_01834_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07527_ (.A1(_01818_),
    .A2(_01834_),
    .ZN(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07528_ (.I(_01677_),
    .Z(_01836_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07529_ (.I(_01510_),
    .Z(_01837_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07530_ (.I(_01503_),
    .Z(_01838_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07531_ (.I0(\mod.u_cpu.rf_ram.memory[324][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[325][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[326][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[327][0] ),
    .S0(_01837_),
    .S1(_01838_),
    .Z(_01839_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07532_ (.I0(\mod.u_cpu.rf_ram.memory[340][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[341][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[342][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[343][0] ),
    .S0(_01826_),
    .S1(_01828_),
    .Z(_01840_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07533_ (.I(_01710_),
    .Z(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07534_ (.I0(\mod.u_cpu.rf_ram.memory[320][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[321][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[322][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[323][0] ),
    .S0(_01841_),
    .S1(_01763_),
    .Z(_01842_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07535_ (.I(_01825_),
    .Z(_01843_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07536_ (.I(_01503_),
    .Z(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07537_ (.I0(\mod.u_cpu.rf_ram.memory[336][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[337][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[338][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[339][0] ),
    .S0(_01843_),
    .S1(_01844_),
    .Z(_01845_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07538_ (.I0(_01839_),
    .I1(_01840_),
    .I2(_01842_),
    .I3(_01845_),
    .S0(_01832_),
    .S1(_01833_),
    .Z(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07539_ (.A1(_01836_),
    .A2(_01846_),
    .B(_01485_),
    .ZN(_01847_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07540_ (.I(_01457_),
    .Z(_01848_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07541_ (.I(_01832_),
    .Z(_01849_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07542_ (.I(_01490_),
    .Z(_01850_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07543_ (.I(_01850_),
    .Z(_01851_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07544_ (.I(_01851_),
    .Z(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07545_ (.I0(\mod.u_cpu.rf_ram.memory[376][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[377][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[378][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[379][0] ),
    .S0(_01837_),
    .S1(_01838_),
    .Z(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07546_ (.I(_01499_),
    .Z(_01854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07547_ (.I(_01854_),
    .Z(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07548_ (.I(_01603_),
    .Z(_01856_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07549_ (.I(_01856_),
    .Z(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07550_ (.I(_01758_),
    .Z(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07551_ (.I(\mod.u_cpu.rf_ram.memory[381][0] ),
    .ZN(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07552_ (.A1(_01858_),
    .A2(_01859_),
    .ZN(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07553_ (.A1(_01857_),
    .A2(\mod.u_cpu.rf_ram.memory[380][0] ),
    .B(_01860_),
    .ZN(_01861_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07554_ (.I(_01509_),
    .Z(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07555_ (.I(_01862_),
    .Z(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07556_ (.I(_01671_),
    .Z(_01864_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07557_ (.I(\mod.u_cpu.rf_ram.memory[383][0] ),
    .ZN(_01865_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07558_ (.A1(_01864_),
    .A2(_01865_),
    .ZN(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07559_ (.I(_01503_),
    .Z(_01867_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07560_ (.A1(_01863_),
    .A2(\mod.u_cpu.rf_ram.memory[382][0] ),
    .B(_01866_),
    .C(_01867_),
    .ZN(_01868_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07561_ (.A1(_01855_),
    .A2(_01861_),
    .B(_01868_),
    .C(_01631_),
    .ZN(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07562_ (.I(_01550_),
    .Z(_01870_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07563_ (.A1(_01852_),
    .A2(_01853_),
    .B(_01869_),
    .C(_01870_),
    .ZN(_01871_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07564_ (.I(_01851_),
    .Z(_01872_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07565_ (.I0(\mod.u_cpu.rf_ram.memory[368][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[369][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[370][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[371][0] ),
    .S0(_01843_),
    .S1(_01844_),
    .Z(_01873_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07566_ (.I(_01665_),
    .Z(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07567_ (.I(_01825_),
    .Z(_01875_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07568_ (.I(\mod.u_cpu.rf_ram.memory[373][0] ),
    .ZN(_01876_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07569_ (.A1(_01759_),
    .A2(_01876_),
    .ZN(_01877_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07570_ (.A1(_01875_),
    .A2(\mod.u_cpu.rf_ram.memory[372][0] ),
    .B(_01877_),
    .ZN(_01878_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07571_ (.I(_01710_),
    .Z(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07572_ (.I(\mod.u_cpu.rf_ram.memory[375][0] ),
    .ZN(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07573_ (.A1(_01663_),
    .A2(_01880_),
    .ZN(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07574_ (.I(_01749_),
    .Z(_01882_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07575_ (.A1(_01879_),
    .A2(\mod.u_cpu.rf_ram.memory[374][0] ),
    .B(_01881_),
    .C(_01882_),
    .ZN(_01883_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07576_ (.I(_01630_),
    .Z(_01884_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07577_ (.A1(_01874_),
    .A2(_01878_),
    .B(_01883_),
    .C(_01884_),
    .ZN(_01885_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07578_ (.I(_01532_),
    .Z(_01886_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07579_ (.I(_01886_),
    .Z(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07580_ (.A1(_01872_),
    .A2(_01873_),
    .B(_01885_),
    .C(_01887_),
    .ZN(_01888_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07581_ (.A1(_01849_),
    .A2(_01871_),
    .A3(_01888_),
    .ZN(_01889_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07582_ (.I(_01487_),
    .Z(_01890_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07583_ (.I(_01890_),
    .Z(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07584_ (.I0(\mod.u_cpu.rf_ram.memory[360][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[361][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[362][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[363][0] ),
    .S0(_01843_),
    .S1(_01838_),
    .Z(_01892_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07585_ (.I(_01856_),
    .Z(_01893_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07586_ (.I(\mod.u_cpu.rf_ram.memory[365][0] ),
    .ZN(_01894_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07587_ (.A1(_01759_),
    .A2(_01894_),
    .ZN(_01895_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07588_ (.A1(_01893_),
    .A2(\mod.u_cpu.rf_ram.memory[364][0] ),
    .B(_01895_),
    .ZN(_01896_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07589_ (.I(\mod.u_cpu.rf_ram.memory[367][0] ),
    .ZN(_01897_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07590_ (.A1(_01663_),
    .A2(_01897_),
    .ZN(_01898_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07591_ (.A1(_01879_),
    .A2(\mod.u_cpu.rf_ram.memory[366][0] ),
    .B(_01898_),
    .C(_01867_),
    .ZN(_01899_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07592_ (.A1(_01874_),
    .A2(_01896_),
    .B(_01899_),
    .C(_01884_),
    .ZN(_01900_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07593_ (.A1(_01852_),
    .A2(_01892_),
    .B(_01900_),
    .C(_01677_),
    .ZN(_01901_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07594_ (.I0(\mod.u_cpu.rf_ram.memory[352][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[353][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[354][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[355][0] ),
    .S0(_01841_),
    .S1(_01844_),
    .Z(_01902_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07595_ (.I(\mod.u_cpu.rf_ram.memory[357][0] ),
    .ZN(_01903_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07596_ (.A1(_01759_),
    .A2(_01903_),
    .ZN(_01904_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07597_ (.A1(_01875_),
    .A2(\mod.u_cpu.rf_ram.memory[356][0] ),
    .B(_01904_),
    .ZN(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07598_ (.I(\mod.u_cpu.rf_ram.memory[359][0] ),
    .ZN(_01906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07599_ (.A1(_01663_),
    .A2(_01906_),
    .ZN(_01907_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07600_ (.A1(_01745_),
    .A2(\mod.u_cpu.rf_ram.memory[358][0] ),
    .B(_01907_),
    .C(_01882_),
    .ZN(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07601_ (.A1(_01874_),
    .A2(_01905_),
    .B(_01908_),
    .C(_01884_),
    .ZN(_01909_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07602_ (.A1(_01872_),
    .A2(_01902_),
    .B(_01909_),
    .C(_01657_),
    .ZN(_01910_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07603_ (.A1(_01891_),
    .A2(_01901_),
    .A3(_01910_),
    .ZN(_01911_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07604_ (.A1(_01848_),
    .A2(_01889_),
    .A3(_01911_),
    .ZN(_01912_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07605_ (.A1(_01835_),
    .A2(_01847_),
    .B(_01912_),
    .C(_01482_),
    .ZN(_01913_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07606_ (.I(_01850_),
    .Z(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07607_ (.I(_01914_),
    .Z(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07608_ (.I(_01581_),
    .Z(_01916_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07609_ (.I0(\mod.u_cpu.rf_ram.memory[312][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[313][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[314][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[315][0] ),
    .S0(_01774_),
    .S1(_01916_),
    .Z(_01917_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07610_ (.I(_01750_),
    .Z(_01918_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07611_ (.I(_01743_),
    .Z(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07612_ (.I(_01919_),
    .Z(_01920_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07613_ (.I(\mod.u_cpu.rf_ram.memory[317][0] ),
    .ZN(_01921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07614_ (.A1(_01920_),
    .A2(_01921_),
    .ZN(_01922_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07615_ (.A1(_01643_),
    .A2(\mod.u_cpu.rf_ram.memory[316][0] ),
    .B(_01922_),
    .ZN(_01923_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07616_ (.I(_01634_),
    .Z(_01924_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07617_ (.I(_01924_),
    .Z(_01925_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07618_ (.I(\mod.u_cpu.rf_ram.memory[319][0] ),
    .ZN(_01926_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07619_ (.A1(_01507_),
    .A2(_01926_),
    .ZN(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07620_ (.A1(_01925_),
    .A2(\mod.u_cpu.rf_ram.memory[318][0] ),
    .B(_01927_),
    .C(_01783_),
    .ZN(_01928_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07621_ (.I(_01686_),
    .Z(_01929_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07622_ (.A1(_01918_),
    .A2(_01923_),
    .B(_01928_),
    .C(_01929_),
    .ZN(_01930_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07623_ (.A1(_01915_),
    .A2(_01917_),
    .B(_01930_),
    .C(_01812_),
    .ZN(_01931_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07624_ (.I(_01827_),
    .Z(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07625_ (.I0(\mod.u_cpu.rf_ram.memory[304][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[305][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[306][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[307][0] ),
    .S0(_01802_),
    .S1(_01932_),
    .Z(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07626_ (.I(_01710_),
    .Z(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07627_ (.I(\mod.u_cpu.rf_ram.memory[309][0] ),
    .ZN(_01935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07628_ (.A1(_01934_),
    .A2(_01935_),
    .ZN(_01936_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07629_ (.A1(_01643_),
    .A2(\mod.u_cpu.rf_ram.memory[308][0] ),
    .B(_01936_),
    .ZN(_01937_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07630_ (.I(_01825_),
    .Z(_01938_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07631_ (.I(\mod.u_cpu.rf_ram.memory[311][0] ),
    .ZN(_01939_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07632_ (.A1(_01507_),
    .A2(_01939_),
    .ZN(_01940_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07633_ (.A1(_01938_),
    .A2(\mod.u_cpu.rf_ram.memory[310][0] ),
    .B(_01940_),
    .C(_01783_),
    .ZN(_01941_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07634_ (.A1(_01918_),
    .A2(_01937_),
    .B(_01941_),
    .C(_01929_),
    .ZN(_01942_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07635_ (.A1(_01915_),
    .A2(_01933_),
    .B(_01942_),
    .C(_01768_),
    .ZN(_01943_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07636_ (.A1(_01791_),
    .A2(_01931_),
    .A3(_01943_),
    .ZN(_01944_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07637_ (.I0(\mod.u_cpu.rf_ram.memory[288][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[289][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[290][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[291][0] ),
    .S0(_01774_),
    .S1(_01932_),
    .Z(_01945_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07638_ (.I(\mod.u_cpu.rf_ram.memory[293][0] ),
    .ZN(_01946_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07639_ (.A1(_01934_),
    .A2(_01946_),
    .ZN(_01947_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07640_ (.A1(_01643_),
    .A2(\mod.u_cpu.rf_ram.memory[292][0] ),
    .B(_01947_),
    .ZN(_01948_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07641_ (.I(_01758_),
    .Z(_01949_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07642_ (.I(\mod.u_cpu.rf_ram.memory[295][0] ),
    .ZN(_01950_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07643_ (.A1(_01949_),
    .A2(_01950_),
    .ZN(_01951_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07644_ (.I(_01782_),
    .Z(_01952_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07645_ (.A1(_01938_),
    .A2(\mod.u_cpu.rf_ram.memory[294][0] ),
    .B(_01951_),
    .C(_01952_),
    .ZN(_01953_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07646_ (.A1(_01918_),
    .A2(_01948_),
    .B(_01953_),
    .C(_01929_),
    .ZN(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07647_ (.A1(_01915_),
    .A2(_01945_),
    .B(_01954_),
    .C(_01768_),
    .ZN(_01955_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07648_ (.I(_01914_),
    .Z(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07649_ (.I(_01919_),
    .Z(_01957_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07650_ (.I(_01827_),
    .Z(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07651_ (.I0(\mod.u_cpu.rf_ram.memory[296][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[297][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[298][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[299][0] ),
    .S0(_01957_),
    .S1(_01958_),
    .Z(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07652_ (.I(_01749_),
    .Z(_01960_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07653_ (.I(_01960_),
    .Z(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07654_ (.I(_01752_),
    .Z(_01962_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07655_ (.I(_01644_),
    .Z(_01963_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07656_ (.I(\mod.u_cpu.rf_ram.memory[301][0] ),
    .ZN(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07657_ (.A1(_01963_),
    .A2(_01964_),
    .ZN(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07658_ (.A1(_01962_),
    .A2(\mod.u_cpu.rf_ram.memory[300][0] ),
    .B(_01965_),
    .ZN(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07659_ (.I(_01758_),
    .Z(_01967_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07660_ (.I(\mod.u_cpu.rf_ram.memory[303][0] ),
    .ZN(_01968_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07661_ (.A1(_01967_),
    .A2(_01968_),
    .ZN(_01969_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07662_ (.I(_01701_),
    .Z(_01970_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07663_ (.A1(_01697_),
    .A2(\mod.u_cpu.rf_ram.memory[302][0] ),
    .B(_01969_),
    .C(_01970_),
    .ZN(_01971_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07664_ (.I(_01686_),
    .Z(_01972_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07665_ (.A1(_01961_),
    .A2(_01966_),
    .B(_01971_),
    .C(_01972_),
    .ZN(_01973_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07666_ (.A1(_01956_),
    .A2(_01959_),
    .B(_01973_),
    .C(_01812_),
    .ZN(_01974_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07667_ (.A1(_01740_),
    .A2(_01955_),
    .A3(_01974_),
    .ZN(_01975_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07668_ (.A1(_01739_),
    .A2(_01944_),
    .A3(_01975_),
    .ZN(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07669_ (.I(_01484_),
    .Z(_01977_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07670_ (.I(_01832_),
    .Z(_01978_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07671_ (.I(_01914_),
    .Z(_01979_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07672_ (.I0(\mod.u_cpu.rf_ram.memory[272][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[273][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[274][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[275][0] ),
    .S0(_01957_),
    .S1(_01958_),
    .Z(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07673_ (.I(_01750_),
    .Z(_01981_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07674_ (.I(\mod.u_cpu.rf_ram.memory[277][0] ),
    .ZN(_01982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07675_ (.A1(_01934_),
    .A2(_01982_),
    .ZN(_01983_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07676_ (.A1(_01962_),
    .A2(\mod.u_cpu.rf_ram.memory[276][0] ),
    .B(_01983_),
    .ZN(_01984_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07677_ (.I(\mod.u_cpu.rf_ram.memory[279][0] ),
    .ZN(_01985_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07678_ (.A1(_01949_),
    .A2(_01985_),
    .ZN(_01986_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07679_ (.A1(_01938_),
    .A2(\mod.u_cpu.rf_ram.memory[278][0] ),
    .B(_01986_),
    .C(_01952_),
    .ZN(_01987_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07680_ (.A1(_01981_),
    .A2(_01984_),
    .B(_01987_),
    .C(_01972_),
    .ZN(_01988_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07681_ (.I(_01886_),
    .Z(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07682_ (.A1(_01979_),
    .A2(_01980_),
    .B(_01988_),
    .C(_01989_),
    .ZN(_01990_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07683_ (.I(_01850_),
    .Z(_01991_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07684_ (.I(_01991_),
    .Z(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07685_ (.I(_01645_),
    .Z(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07686_ (.I(_01993_),
    .Z(_01994_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07687_ (.I(_01762_),
    .Z(_01995_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07688_ (.I0(\mod.u_cpu.rf_ram.memory[280][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[281][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[282][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[283][0] ),
    .S0(_01994_),
    .S1(_01995_),
    .Z(_01996_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07689_ (.I(_01960_),
    .Z(_01997_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07690_ (.I(_01752_),
    .Z(_01998_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07691_ (.I(\mod.u_cpu.rf_ram.memory[285][0] ),
    .ZN(_01999_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07692_ (.A1(_01711_),
    .A2(_01999_),
    .ZN(_02000_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07693_ (.A1(_01998_),
    .A2(\mod.u_cpu.rf_ram.memory[284][0] ),
    .B(_02000_),
    .ZN(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07694_ (.I(\mod.u_cpu.rf_ram.memory[287][0] ),
    .ZN(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07695_ (.A1(_01967_),
    .A2(_02002_),
    .ZN(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07696_ (.A1(_01722_),
    .A2(\mod.u_cpu.rf_ram.memory[286][0] ),
    .B(_02003_),
    .C(_01970_),
    .ZN(_02004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07697_ (.I(_01491_),
    .Z(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07698_ (.A1(_01997_),
    .A2(_02001_),
    .B(_02004_),
    .C(_02005_),
    .ZN(_02006_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07699_ (.I(_01787_),
    .Z(_02007_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07700_ (.A1(_01992_),
    .A2(_01996_),
    .B(_02006_),
    .C(_02007_),
    .ZN(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07701_ (.A1(_01978_),
    .A2(_01990_),
    .A3(_02008_),
    .ZN(_02009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07702_ (.I(_01581_),
    .Z(_02010_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07703_ (.I0(\mod.u_cpu.rf_ram.memory[256][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[257][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[258][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[259][0] ),
    .S0(_01994_),
    .S1(_02010_),
    .Z(_02011_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07704_ (.I(\mod.u_cpu.rf_ram.memory[261][0] ),
    .ZN(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07705_ (.A1(_01711_),
    .A2(_02012_),
    .ZN(_02013_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07706_ (.A1(_01998_),
    .A2(\mod.u_cpu.rf_ram.memory[260][0] ),
    .B(_02013_),
    .ZN(_02014_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07707_ (.I(\mod.u_cpu.rf_ram.memory[263][0] ),
    .ZN(_02015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07708_ (.A1(_01967_),
    .A2(_02015_),
    .ZN(_02016_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07709_ (.A1(_01722_),
    .A2(\mod.u_cpu.rf_ram.memory[262][0] ),
    .B(_02016_),
    .C(_01970_),
    .ZN(_02017_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07710_ (.A1(_01961_),
    .A2(_02014_),
    .B(_02017_),
    .C(_02005_),
    .ZN(_02018_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07711_ (.A1(_01956_),
    .A2(_02011_),
    .B(_02018_),
    .C(_01989_),
    .ZN(_02019_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07712_ (.I(_01993_),
    .Z(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07713_ (.I0(\mod.u_cpu.rf_ram.memory[264][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[265][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[266][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[267][0] ),
    .S0(_02020_),
    .S1(_01995_),
    .Z(_02021_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07714_ (.I(_01704_),
    .Z(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07715_ (.I(\mod.u_cpu.rf_ram.memory[269][0] ),
    .ZN(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07716_ (.A1(_01729_),
    .A2(_02023_),
    .ZN(_02024_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07717_ (.A1(_02022_),
    .A2(\mod.u_cpu.rf_ram.memory[268][0] ),
    .B(_02024_),
    .ZN(_02025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07718_ (.I(_01757_),
    .Z(_02026_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07719_ (.I(_02026_),
    .Z(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07720_ (.I(\mod.u_cpu.rf_ram.memory[271][0] ),
    .ZN(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07721_ (.A1(_02027_),
    .A2(_02028_),
    .ZN(_02029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07722_ (.I(_01782_),
    .Z(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07723_ (.A1(_01857_),
    .A2(\mod.u_cpu.rf_ram.memory[270][0] ),
    .B(_02029_),
    .C(_02030_),
    .ZN(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07724_ (.A1(_01997_),
    .A2(_02025_),
    .B(_02031_),
    .C(_02005_),
    .ZN(_02032_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07725_ (.A1(_01992_),
    .A2(_02021_),
    .B(_02032_),
    .C(_02007_),
    .ZN(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07726_ (.A1(_01740_),
    .A2(_02019_),
    .A3(_02033_),
    .ZN(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07727_ (.A1(_01977_),
    .A2(_02009_),
    .A3(_02034_),
    .ZN(_02035_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07728_ (.A1(_01738_),
    .A2(_01976_),
    .A3(_02035_),
    .ZN(_02036_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07729_ (.A1(_01471_),
    .A2(_01913_),
    .A3(_02036_),
    .Z(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07730_ (.A1(_01481_),
    .A2(_01817_),
    .B(_02037_),
    .C(_01469_),
    .ZN(_02038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07731_ (.I(_01485_),
    .Z(_02039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07732_ (.I(_01444_),
    .Z(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07733_ (.I(_01743_),
    .Z(_02041_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07734_ (.I(_01499_),
    .Z(_02042_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07735_ (.I(_02042_),
    .Z(_02043_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07736_ (.I0(\mod.u_cpu.rf_ram.memory[128][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[129][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[130][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[131][0] ),
    .S0(_02041_),
    .S1(_02043_),
    .Z(_02044_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07737_ (.A1(_02040_),
    .A2(_02044_),
    .ZN(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07738_ (.I(_01890_),
    .Z(_02046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07739_ (.I(_02026_),
    .Z(_02047_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07740_ (.I(_02047_),
    .Z(_02048_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07741_ (.I(_02042_),
    .Z(_02049_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07742_ (.I0(\mod.u_cpu.rf_ram.memory[144][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[145][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[146][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[147][0] ),
    .S0(_02048_),
    .S1(_02049_),
    .Z(_02050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07743_ (.I(_01661_),
    .Z(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07744_ (.A1(_02046_),
    .A2(_02050_),
    .B(_02051_),
    .ZN(_02052_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07745_ (.I(_01444_),
    .Z(_02053_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07746_ (.I(_01569_),
    .Z(_02054_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07747_ (.I0(\mod.u_cpu.rf_ram.memory[132][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[133][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[134][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[135][0] ),
    .S0(_01893_),
    .S1(_02054_),
    .Z(_02055_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07748_ (.A1(_02053_),
    .A2(_02055_),
    .ZN(_02056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07749_ (.I(_01487_),
    .Z(_02057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07750_ (.I(_01603_),
    .Z(_02058_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07751_ (.I(_02058_),
    .Z(_02059_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07752_ (.I0(\mod.u_cpu.rf_ram.memory[148][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[149][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[150][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[151][0] ),
    .S0(_02059_),
    .S1(_01723_),
    .Z(_02060_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07753_ (.A1(_02057_),
    .A2(_02060_),
    .B(_01632_),
    .ZN(_02061_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07754_ (.A1(_02045_),
    .A2(_02052_),
    .B1(_02056_),
    .B2(_02061_),
    .C(_01818_),
    .ZN(_02062_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07755_ (.I(_01960_),
    .Z(_02063_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07756_ (.I0(\mod.u_cpu.rf_ram.memory[136][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[137][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[138][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[139][0] ),
    .S0(_02022_),
    .S1(_02063_),
    .Z(_02064_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07757_ (.A1(_01849_),
    .A2(_02064_),
    .ZN(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07758_ (.I(_01704_),
    .Z(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07759_ (.I(_02042_),
    .Z(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07760_ (.I0(\mod.u_cpu.rf_ram.memory[152][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[153][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[154][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[155][0] ),
    .S0(_02066_),
    .S1(_02067_),
    .Z(_02068_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07761_ (.A1(_02046_),
    .A2(_02068_),
    .B(_02051_),
    .ZN(_02069_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07762_ (.I(_01806_),
    .Z(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07763_ (.I(_01746_),
    .Z(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07764_ (.I0(\mod.u_cpu.rf_ram.memory[140][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[141][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[142][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[143][0] ),
    .S0(_02070_),
    .S1(_02071_),
    .Z(_02072_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07765_ (.A1(_02053_),
    .A2(_02072_),
    .ZN(_02073_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07766_ (.I(_01890_),
    .Z(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07767_ (.I0(\mod.u_cpu.rf_ram.memory[156][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[157][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[158][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[159][0] ),
    .S0(_01925_),
    .S1(_02071_),
    .Z(_02075_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07768_ (.A1(_02074_),
    .A2(_02075_),
    .B(_01602_),
    .ZN(_02076_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07769_ (.I(_01677_),
    .Z(_02077_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07770_ (.A1(_02065_),
    .A2(_02069_),
    .B1(_02073_),
    .B2(_02076_),
    .C(_02077_),
    .ZN(_02078_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07771_ (.A1(_02039_),
    .A2(_02062_),
    .A3(_02078_),
    .Z(_02079_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07772_ (.I(_01661_),
    .Z(_02080_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07773_ (.I0(\mod.u_cpu.rf_ram.memory[176][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[177][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[178][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[179][0] ),
    .S0(_02048_),
    .S1(_02049_),
    .Z(_02081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07774_ (.A1(_02080_),
    .A2(_02081_),
    .ZN(_02082_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07775_ (.I(_01785_),
    .Z(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07776_ (.I(_01671_),
    .Z(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07777_ (.I(_02084_),
    .Z(_02085_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07778_ (.I(_01854_),
    .Z(_02086_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07779_ (.I0(\mod.u_cpu.rf_ram.memory[180][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[181][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[182][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[183][0] ),
    .S0(_02085_),
    .S1(_02086_),
    .Z(_02087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07780_ (.A1(_02083_),
    .A2(_02087_),
    .ZN(_02088_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07781_ (.A1(_01818_),
    .A2(_02082_),
    .A3(_02088_),
    .ZN(_02089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07782_ (.I(_01661_),
    .Z(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07783_ (.I(_01671_),
    .Z(_02091_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07784_ (.I(_02091_),
    .Z(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07785_ (.I(_02042_),
    .Z(_02093_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07786_ (.I0(\mod.u_cpu.rf_ram.memory[184][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[185][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[186][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[187][0] ),
    .S0(_02092_),
    .S1(_02093_),
    .Z(_02094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07787_ (.A1(_02090_),
    .A2(_02094_),
    .ZN(_02095_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07788_ (.I(_01686_),
    .Z(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07789_ (.I(_02096_),
    .Z(_02097_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07790_ (.I(_01637_),
    .Z(_02098_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07791_ (.I0(\mod.u_cpu.rf_ram.memory[188][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[189][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[190][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[191][0] ),
    .S0(_02092_),
    .S1(_02098_),
    .Z(_02099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07792_ (.A1(_02097_),
    .A2(_02099_),
    .ZN(_02100_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07793_ (.A1(_01836_),
    .A2(_02095_),
    .A3(_02100_),
    .ZN(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07794_ (.I(_02057_),
    .Z(_02102_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07795_ (.A1(_02089_),
    .A2(_02101_),
    .B(_02102_),
    .ZN(_02103_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07796_ (.I(_01458_),
    .Z(_02104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07797_ (.I(_01488_),
    .Z(_02105_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07798_ (.I(_01672_),
    .Z(_02106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07799_ (.I(_01854_),
    .Z(_02107_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07800_ (.I0(\mod.u_cpu.rf_ram.memory[168][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[169][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[170][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[171][0] ),
    .S0(_02106_),
    .S1(_02107_),
    .Z(_02108_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07801_ (.I(_01701_),
    .Z(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07802_ (.I(_02109_),
    .Z(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07803_ (.I(_02047_),
    .Z(_02111_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07804_ (.I(\mod.u_cpu.rf_ram.memory[173][0] ),
    .ZN(_02112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07805_ (.A1(_01673_),
    .A2(_02112_),
    .ZN(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07806_ (.A1(_02111_),
    .A2(\mod.u_cpu.rf_ram.memory[172][0] ),
    .B(_02113_),
    .ZN(_02114_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07807_ (.I(_01635_),
    .Z(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07808_ (.I(_01862_),
    .Z(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07809_ (.I(\mod.u_cpu.rf_ram.memory[175][0] ),
    .ZN(_02117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07810_ (.A1(_02116_),
    .A2(_02117_),
    .ZN(_02118_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07811_ (.A1(_02115_),
    .A2(\mod.u_cpu.rf_ram.memory[174][0] ),
    .B(_02118_),
    .C(_01771_),
    .ZN(_02119_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07812_ (.I(_01716_),
    .Z(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07813_ (.A1(_02110_),
    .A2(_02114_),
    .B(_02119_),
    .C(_02120_),
    .ZN(_02121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07814_ (.I(_01719_),
    .Z(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07815_ (.A1(_01670_),
    .A2(_02108_),
    .B(_02121_),
    .C(_02122_),
    .ZN(_02123_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07816_ (.I(_01687_),
    .Z(_02124_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07817_ (.I(_01672_),
    .Z(_02125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07818_ (.I(_01568_),
    .Z(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07819_ (.I(_02126_),
    .Z(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07820_ (.I0(\mod.u_cpu.rf_ram.memory[160][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[161][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[162][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[163][0] ),
    .S0(_02125_),
    .S1(_02127_),
    .Z(_02128_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07821_ (.I(_02047_),
    .Z(_02129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07822_ (.I(_01744_),
    .Z(_02130_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07823_ (.I(\mod.u_cpu.rf_ram.memory[165][0] ),
    .ZN(_02131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07824_ (.A1(_02130_),
    .A2(_02131_),
    .ZN(_02132_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07825_ (.A1(_02129_),
    .A2(\mod.u_cpu.rf_ram.memory[164][0] ),
    .B(_02132_),
    .ZN(_02133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07826_ (.I(_01634_),
    .Z(_02134_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07827_ (.I(_02134_),
    .Z(_02135_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07828_ (.I(_01862_),
    .Z(_02136_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07829_ (.I(\mod.u_cpu.rf_ram.memory[167][0] ),
    .ZN(_02137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07830_ (.A1(_02136_),
    .A2(_02137_),
    .ZN(_02138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07831_ (.I(_01746_),
    .Z(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07832_ (.A1(_02135_),
    .A2(\mod.u_cpu.rf_ram.memory[166][0] ),
    .B(_02138_),
    .C(_02139_),
    .ZN(_02140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07833_ (.I(_01716_),
    .Z(_02141_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07834_ (.A1(_02110_),
    .A2(_02133_),
    .B(_02140_),
    .C(_02141_),
    .ZN(_02142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07835_ (.I(_01533_),
    .Z(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07836_ (.A1(_02124_),
    .A2(_02128_),
    .B(_02142_),
    .C(_02143_),
    .ZN(_02144_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07837_ (.A1(_02105_),
    .A2(_02123_),
    .A3(_02144_),
    .ZN(_02145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07838_ (.A1(_02104_),
    .A2(_02145_),
    .ZN(_02146_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07839_ (.A1(_02103_),
    .A2(_02146_),
    .B(_01475_),
    .ZN(_02147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07840_ (.I(_01482_),
    .Z(_02148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07841_ (.I(_01488_),
    .Z(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07842_ (.I(_01741_),
    .Z(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07843_ (.I(_01856_),
    .Z(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07844_ (.I(_02126_),
    .Z(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07845_ (.I0(\mod.u_cpu.rf_ram.memory[192][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[193][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[194][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[195][0] ),
    .S0(_02151_),
    .S1(_02152_),
    .Z(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07846_ (.I(_01749_),
    .Z(_02154_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07847_ (.I(_02154_),
    .Z(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07848_ (.I(_01635_),
    .Z(_02156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07849_ (.I(_01681_),
    .Z(_02157_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07850_ (.I(\mod.u_cpu.rf_ram.memory[197][0] ),
    .ZN(_02158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07851_ (.A1(_02157_),
    .A2(_02158_),
    .ZN(_02159_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07852_ (.A1(_02156_),
    .A2(\mod.u_cpu.rf_ram.memory[196][0] ),
    .B(_02159_),
    .ZN(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07853_ (.I(_01646_),
    .Z(_02161_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07854_ (.I(\mod.u_cpu.rf_ram.memory[199][0] ),
    .ZN(_02162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07855_ (.A1(_01819_),
    .A2(_02162_),
    .ZN(_02163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07856_ (.I(_01820_),
    .Z(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07857_ (.A1(_02161_),
    .A2(\mod.u_cpu.rf_ram.memory[198][0] ),
    .B(_02163_),
    .C(_02164_),
    .ZN(_02165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07858_ (.I(_01765_),
    .Z(_02166_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07859_ (.A1(_02155_),
    .A2(_02160_),
    .B(_02165_),
    .C(_02166_),
    .ZN(_02167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07860_ (.I(_01586_),
    .Z(_02168_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07861_ (.A1(_02150_),
    .A2(_02153_),
    .B(_02167_),
    .C(_02168_),
    .ZN(_02169_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07862_ (.I(_01741_),
    .Z(_02170_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07863_ (.I(_01806_),
    .Z(_02171_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07864_ (.I(_01614_),
    .Z(_02172_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07865_ (.I0(\mod.u_cpu.rf_ram.memory[200][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[201][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[202][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[203][0] ),
    .S0(_02171_),
    .S1(_02172_),
    .Z(_02173_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07866_ (.I(_02154_),
    .Z(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07867_ (.I(_02134_),
    .Z(_02175_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07868_ (.I(\mod.u_cpu.rf_ram.memory[205][0] ),
    .ZN(_02176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07869_ (.A1(_02157_),
    .A2(_02176_),
    .ZN(_02177_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07870_ (.A1(_02175_),
    .A2(\mod.u_cpu.rf_ram.memory[204][0] ),
    .B(_02177_),
    .ZN(_02178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07871_ (.I(_01646_),
    .Z(_02179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07872_ (.I(_01778_),
    .Z(_02180_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07873_ (.I(\mod.u_cpu.rf_ram.memory[207][0] ),
    .ZN(_02181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07874_ (.A1(_02180_),
    .A2(_02181_),
    .ZN(_02182_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07875_ (.A1(_02179_),
    .A2(\mod.u_cpu.rf_ram.memory[206][0] ),
    .B(_02182_),
    .C(_02164_),
    .ZN(_02183_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07876_ (.A1(_02174_),
    .A2(_02178_),
    .B(_02183_),
    .C(_02166_),
    .ZN(_02184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07877_ (.I(_01551_),
    .Z(_02185_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07878_ (.A1(_02170_),
    .A2(_02173_),
    .B(_02184_),
    .C(_02185_),
    .ZN(_02186_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07879_ (.A1(_02149_),
    .A2(_02169_),
    .A3(_02186_),
    .ZN(_02187_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07880_ (.I(_01582_),
    .Z(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07881_ (.I0(\mod.u_cpu.rf_ram.memory[222][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[223][0] ),
    .S(_02048_),
    .Z(_02189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07882_ (.I(_02026_),
    .Z(_02190_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07883_ (.I(_02190_),
    .Z(_02191_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07884_ (.I(\mod.u_cpu.rf_ram.memory[221][0] ),
    .ZN(_02192_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07885_ (.A1(_01682_),
    .A2(\mod.u_cpu.rf_ram.memory[220][0] ),
    .ZN(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07886_ (.A1(_02191_),
    .A2(_02192_),
    .B(_02193_),
    .C(_01666_),
    .ZN(_02194_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07887_ (.A1(_02188_),
    .A2(_02189_),
    .B(_02194_),
    .C(_01833_),
    .ZN(_02195_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07888_ (.I(_01851_),
    .Z(_02196_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07889_ (.I(_01519_),
    .Z(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07890_ (.I(_02197_),
    .Z(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07891_ (.I(\mod.u_cpu.rf_ram.memory[219][0] ),
    .ZN(_02199_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07892_ (.A1(_01517_),
    .A2(\mod.u_cpu.rf_ram.memory[218][0] ),
    .B(_01714_),
    .ZN(_02200_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07893_ (.A1(_02198_),
    .A2(_02199_),
    .B(_02200_),
    .ZN(_02201_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07894_ (.I(_01779_),
    .Z(_02202_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07895_ (.I(\mod.u_cpu.rf_ram.memory[217][0] ),
    .ZN(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07896_ (.I(_01993_),
    .Z(_02204_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07897_ (.A1(_02204_),
    .A2(\mod.u_cpu.rf_ram.memory[216][0] ),
    .ZN(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07898_ (.A1(_02202_),
    .A2(_02203_),
    .B(_02205_),
    .C(_02049_),
    .ZN(_02206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07899_ (.I(_01787_),
    .Z(_02207_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _07900_ (.A1(_02196_),
    .A2(_02201_),
    .A3(_02206_),
    .B(_02207_),
    .ZN(_02208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07901_ (.I(_02091_),
    .Z(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07902_ (.I(\mod.u_cpu.rf_ram.memory[211][0] ),
    .ZN(_02210_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07903_ (.I(_01924_),
    .Z(_02211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07904_ (.I(_01701_),
    .Z(_02212_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07905_ (.A1(_02211_),
    .A2(\mod.u_cpu.rf_ram.memory[210][0] ),
    .B(_02212_),
    .ZN(_02213_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07906_ (.A1(_02209_),
    .A2(_02210_),
    .B(_02213_),
    .ZN(_02214_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07907_ (.I(\mod.u_cpu.rf_ram.memory[209][0] ),
    .ZN(_02215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07908_ (.I(_01681_),
    .Z(_02216_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07909_ (.A1(_02216_),
    .A2(\mod.u_cpu.rf_ram.memory[208][0] ),
    .ZN(_02217_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07910_ (.I(_01746_),
    .Z(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07911_ (.A1(_01607_),
    .A2(_02215_),
    .B(_02217_),
    .C(_02218_),
    .ZN(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07912_ (.I(_01519_),
    .Z(_02220_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07913_ (.I(\mod.u_cpu.rf_ram.memory[215][0] ),
    .ZN(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07914_ (.A1(_02220_),
    .A2(_02221_),
    .ZN(_02222_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07915_ (.A1(_02066_),
    .A2(\mod.u_cpu.rf_ram.memory[214][0] ),
    .B(_02222_),
    .C(_01821_),
    .ZN(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07916_ (.A1(_01651_),
    .A2(_02223_),
    .ZN(_02224_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07917_ (.I(_01518_),
    .Z(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07918_ (.I(\mod.u_cpu.rf_ram.memory[213][0] ),
    .ZN(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07919_ (.A1(_02070_),
    .A2(\mod.u_cpu.rf_ram.memory[212][0] ),
    .ZN(_02227_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07920_ (.A1(_02225_),
    .A2(_02226_),
    .B(_02227_),
    .C(_01683_),
    .ZN(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _07921_ (.A1(_02120_),
    .A2(_02214_),
    .A3(_02219_),
    .B1(_02224_),
    .B2(_02228_),
    .ZN(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07922_ (.I(_01719_),
    .Z(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07923_ (.A1(_02195_),
    .A2(_02208_),
    .B1(_02229_),
    .B2(_02230_),
    .C(_01978_),
    .ZN(_02231_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07924_ (.A1(_01977_),
    .A2(_02187_),
    .A3(_02231_),
    .ZN(_02232_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07925_ (.I0(\mod.u_cpu.rf_ram.memory[224][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[225][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[226][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[227][0] ),
    .S0(_02151_),
    .S1(_02172_),
    .Z(_02233_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07926_ (.I(\mod.u_cpu.rf_ram.memory[229][0] ),
    .ZN(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07927_ (.A1(_02157_),
    .A2(_02234_),
    .ZN(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07928_ (.A1(_02175_),
    .A2(\mod.u_cpu.rf_ram.memory[228][0] ),
    .B(_02235_),
    .ZN(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07929_ (.I(\mod.u_cpu.rf_ram.memory[231][0] ),
    .ZN(_02237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07930_ (.A1(_01819_),
    .A2(_02237_),
    .ZN(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07931_ (.A1(_02179_),
    .A2(\mod.u_cpu.rf_ram.memory[230][0] ),
    .B(_02238_),
    .C(_02164_),
    .ZN(_02239_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07932_ (.A1(_02155_),
    .A2(_02236_),
    .B(_02239_),
    .C(_02166_),
    .ZN(_02240_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07933_ (.A1(_02170_),
    .A2(_02233_),
    .B(_02240_),
    .C(_02168_),
    .ZN(_02241_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07934_ (.I(_01604_),
    .Z(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07935_ (.I0(\mod.u_cpu.rf_ram.memory[232][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[233][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[234][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[235][0] ),
    .S0(_02242_),
    .S1(_02172_),
    .Z(_02243_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07936_ (.I(_01806_),
    .Z(_02244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07937_ (.I(_01681_),
    .Z(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07938_ (.I(\mod.u_cpu.rf_ram.memory[237][0] ),
    .ZN(_02246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07939_ (.A1(_02245_),
    .A2(_02246_),
    .ZN(_02247_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07940_ (.A1(_02244_),
    .A2(\mod.u_cpu.rf_ram.memory[236][0] ),
    .B(_02247_),
    .ZN(_02248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07941_ (.I(_01539_),
    .Z(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07942_ (.I(\mod.u_cpu.rf_ram.memory[239][0] ),
    .ZN(_02250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07943_ (.A1(_02180_),
    .A2(_02250_),
    .ZN(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07944_ (.I(_01827_),
    .Z(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07945_ (.A1(_02249_),
    .A2(\mod.u_cpu.rf_ram.memory[238][0] ),
    .B(_02251_),
    .C(_02252_),
    .ZN(_02253_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07946_ (.A1(_02174_),
    .A2(_02248_),
    .B(_02253_),
    .C(_01766_),
    .ZN(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07947_ (.A1(_02170_),
    .A2(_02243_),
    .B(_02254_),
    .C(_02207_),
    .ZN(_02255_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07948_ (.A1(_01740_),
    .A2(_02241_),
    .A3(_02255_),
    .ZN(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07949_ (.I0(\mod.u_cpu.rf_ram.memory[240][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[241][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[242][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[243][0] ),
    .S0(_02242_),
    .S1(_02172_),
    .Z(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07950_ (.I(\mod.u_cpu.rf_ram.memory[245][0] ),
    .ZN(_02258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07951_ (.A1(_02245_),
    .A2(_02258_),
    .ZN(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07952_ (.A1(_02175_),
    .A2(\mod.u_cpu.rf_ram.memory[244][0] ),
    .B(_02259_),
    .ZN(_02260_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07953_ (.I(\mod.u_cpu.rf_ram.memory[247][0] ),
    .ZN(_02261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07954_ (.A1(_02180_),
    .A2(_02261_),
    .ZN(_02262_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07955_ (.A1(_02249_),
    .A2(\mod.u_cpu.rf_ram.memory[246][0] ),
    .B(_02262_),
    .C(_02252_),
    .ZN(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07956_ (.A1(_02174_),
    .A2(_02260_),
    .B(_02263_),
    .C(_01766_),
    .ZN(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07957_ (.A1(_02170_),
    .A2(_02257_),
    .B(_02264_),
    .C(_02168_),
    .ZN(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07958_ (.I(_02058_),
    .Z(_02266_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07959_ (.I(_01614_),
    .Z(_02267_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07960_ (.I0(\mod.u_cpu.rf_ram.memory[248][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[249][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[250][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[251][0] ),
    .S0(_02266_),
    .S1(_02267_),
    .Z(_02268_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07961_ (.I(\mod.u_cpu.rf_ram.memory[253][0] ),
    .ZN(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07962_ (.A1(_02245_),
    .A2(_02269_),
    .ZN(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07963_ (.A1(_02244_),
    .A2(\mod.u_cpu.rf_ram.memory[252][0] ),
    .B(_02270_),
    .ZN(_02271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07964_ (.I(_01537_),
    .Z(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07965_ (.I(\mod.u_cpu.rf_ram.memory[255][0] ),
    .ZN(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07966_ (.A1(_02180_),
    .A2(_02273_),
    .ZN(_02274_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07967_ (.A1(_02272_),
    .A2(\mod.u_cpu.rf_ram.memory[254][0] ),
    .B(_02274_),
    .C(_02252_),
    .ZN(_02275_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07968_ (.A1(_02174_),
    .A2(_02271_),
    .B(_02275_),
    .C(_01766_),
    .ZN(_02276_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07969_ (.A1(_01742_),
    .A2(_02268_),
    .B(_02276_),
    .C(_02207_),
    .ZN(_02277_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07970_ (.A1(_01791_),
    .A2(_02265_),
    .A3(_02277_),
    .ZN(_02278_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07971_ (.A1(_01739_),
    .A2(_02256_),
    .A3(_02278_),
    .ZN(_02279_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07972_ (.A1(_02148_),
    .A2(_02232_),
    .A3(_02279_),
    .ZN(_02280_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07973_ (.A1(_02079_),
    .A2(_02147_),
    .B(_01481_),
    .C(_02280_),
    .ZN(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07974_ (.I0(\mod.u_cpu.rf_ram.memory[96][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[97][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[98][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[99][0] ),
    .S0(_02125_),
    .S1(_02127_),
    .Z(_02282_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07975_ (.I(_02212_),
    .Z(_02283_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07976_ (.I(\mod.u_cpu.rf_ram.memory[101][0] ),
    .ZN(_02284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07977_ (.A1(_02130_),
    .A2(_02284_),
    .ZN(_02285_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07978_ (.A1(_02129_),
    .A2(\mod.u_cpu.rf_ram.memory[100][0] ),
    .B(_02285_),
    .ZN(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07979_ (.I(\mod.u_cpu.rf_ram.memory[103][0] ),
    .ZN(_02287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07980_ (.A1(_02136_),
    .A2(_02287_),
    .ZN(_02288_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07981_ (.A1(_02135_),
    .A2(\mod.u_cpu.rf_ram.memory[102][0] ),
    .B(_02288_),
    .C(_02139_),
    .ZN(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07982_ (.A1(_02283_),
    .A2(_02286_),
    .B(_02289_),
    .C(_02141_),
    .ZN(_02290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07983_ (.I(_01533_),
    .Z(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07984_ (.A1(_02124_),
    .A2(_02282_),
    .B(_02290_),
    .C(_02291_),
    .ZN(_02292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07985_ (.I(_01669_),
    .Z(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07986_ (.I(_01864_),
    .Z(_02294_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07987_ (.I(_01854_),
    .Z(_02295_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07988_ (.I0(\mod.u_cpu.rf_ram.memory[104][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[105][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[106][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[107][0] ),
    .S0(_02294_),
    .S1(_02295_),
    .Z(_02296_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07989_ (.I(_02091_),
    .Z(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07990_ (.I(_01744_),
    .Z(_02298_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07991_ (.I(\mod.u_cpu.rf_ram.memory[109][0] ),
    .ZN(_02299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07992_ (.A1(_02298_),
    .A2(_02299_),
    .ZN(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07993_ (.A1(_02297_),
    .A2(\mod.u_cpu.rf_ram.memory[108][0] ),
    .B(_02300_),
    .ZN(_02301_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07994_ (.I(_02134_),
    .Z(_02302_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07995_ (.I(_01862_),
    .Z(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07996_ (.I(\mod.u_cpu.rf_ram.memory[111][0] ),
    .ZN(_02304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07997_ (.A1(_02303_),
    .A2(_02304_),
    .ZN(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07998_ (.I(_01569_),
    .Z(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07999_ (.A1(_02302_),
    .A2(\mod.u_cpu.rf_ram.memory[110][0] ),
    .B(_02305_),
    .C(_02306_),
    .ZN(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08000_ (.I(_01716_),
    .Z(_02308_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08001_ (.A1(_02283_),
    .A2(_02301_),
    .B(_02307_),
    .C(_02308_),
    .ZN(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08002_ (.A1(_02293_),
    .A2(_02296_),
    .B(_02309_),
    .C(_02122_),
    .ZN(_02310_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08003_ (.A1(_02105_),
    .A2(_02292_),
    .A3(_02310_),
    .ZN(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08004_ (.I0(\mod.u_cpu.rf_ram.memory[120][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[121][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[122][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[123][0] ),
    .S0(_02294_),
    .S1(_02295_),
    .Z(_02312_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08005_ (.I(\mod.u_cpu.rf_ram.memory[125][0] ),
    .ZN(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08006_ (.A1(_02298_),
    .A2(_02313_),
    .ZN(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08007_ (.A1(_02297_),
    .A2(\mod.u_cpu.rf_ram.memory[124][0] ),
    .B(_02314_),
    .ZN(_02315_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08008_ (.I(_01924_),
    .Z(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08009_ (.I(\mod.u_cpu.rf_ram.memory[127][0] ),
    .ZN(_02317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08010_ (.A1(_02303_),
    .A2(_02317_),
    .ZN(_02318_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08011_ (.A1(_02316_),
    .A2(\mod.u_cpu.rf_ram.memory[126][0] ),
    .B(_02318_),
    .C(_02306_),
    .ZN(_02319_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08012_ (.A1(_02283_),
    .A2(_02315_),
    .B(_02319_),
    .C(_02308_),
    .ZN(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08013_ (.I(_01719_),
    .Z(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08014_ (.A1(_02293_),
    .A2(_02312_),
    .B(_02320_),
    .C(_02321_),
    .ZN(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08015_ (.I(_01665_),
    .Z(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08016_ (.I0(\mod.u_cpu.rf_ram.memory[112][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[113][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[114][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[115][0] ),
    .S0(_01664_),
    .S1(_02323_),
    .Z(_02324_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08017_ (.I(_02109_),
    .Z(_02325_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08018_ (.I(\mod.u_cpu.rf_ram.memory[117][0] ),
    .ZN(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08019_ (.A1(_02298_),
    .A2(_02326_),
    .ZN(_02327_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08020_ (.A1(_02297_),
    .A2(\mod.u_cpu.rf_ram.memory[116][0] ),
    .B(_02327_),
    .ZN(_02328_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08021_ (.I(_02134_),
    .Z(_02329_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08022_ (.I(\mod.u_cpu.rf_ram.memory[119][0] ),
    .ZN(_02330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08023_ (.A1(_01863_),
    .A2(_02330_),
    .ZN(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08024_ (.A1(_02329_),
    .A2(\mod.u_cpu.rf_ram.memory[118][0] ),
    .B(_02331_),
    .C(_01916_),
    .ZN(_02332_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08025_ (.A1(_02325_),
    .A2(_02328_),
    .B(_02332_),
    .C(_01717_),
    .ZN(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08026_ (.A1(_02293_),
    .A2(_02324_),
    .B(_02333_),
    .C(_02291_),
    .ZN(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08027_ (.A1(_01693_),
    .A2(_02322_),
    .A3(_02334_),
    .ZN(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08028_ (.A1(_02104_),
    .A2(_02311_),
    .A3(_02335_),
    .ZN(_02336_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08029_ (.I(_02057_),
    .Z(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08030_ (.I0(\mod.u_cpu.rf_ram.memory[80][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[81][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[82][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[83][0] ),
    .S0(_02249_),
    .S1(_02098_),
    .Z(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08031_ (.A1(_02090_),
    .A2(_02338_),
    .ZN(_02339_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08032_ (.I0(\mod.u_cpu.rf_ram.memory[84][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[85][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[86][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[87][0] ),
    .S0(_01857_),
    .S1(_02054_),
    .Z(_02340_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08033_ (.A1(_01696_),
    .A2(_02340_),
    .B(_02321_),
    .ZN(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08034_ (.I0(\mod.u_cpu.rf_ram.memory[88][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[89][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[90][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[91][0] ),
    .S0(_01673_),
    .S1(_01666_),
    .Z(_02342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08035_ (.A1(_01662_),
    .A2(_02342_),
    .ZN(_02343_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08036_ (.I0(\mod.u_cpu.rf_ram.memory[92][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[93][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[94][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[95][0] ),
    .S0(_01636_),
    .S1(_01638_),
    .Z(_02344_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08037_ (.A1(_01493_),
    .A2(_02344_),
    .B(_01534_),
    .ZN(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08038_ (.A1(_02339_),
    .A2(_02341_),
    .B1(_02343_),
    .B2(_02345_),
    .ZN(_02346_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08039_ (.I(_01630_),
    .Z(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08040_ (.I(_02347_),
    .Z(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08041_ (.I(_02058_),
    .Z(_02349_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08042_ (.I(_01637_),
    .Z(_02350_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08043_ (.I0(\mod.u_cpu.rf_ram.memory[64][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[65][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[66][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[67][0] ),
    .S0(_02349_),
    .S1(_02350_),
    .Z(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08044_ (.I(_01882_),
    .Z(_02352_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08045_ (.I(\mod.u_cpu.rf_ram.memory[69][0] ),
    .ZN(_02353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08046_ (.A1(_02266_),
    .A2(_02353_),
    .ZN(_02354_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08047_ (.A1(_02135_),
    .A2(\mod.u_cpu.rf_ram.memory[68][0] ),
    .B(_02354_),
    .ZN(_02355_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08048_ (.I(_01993_),
    .Z(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08049_ (.I(\mod.u_cpu.rf_ram.memory[71][0] ),
    .ZN(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08050_ (.A1(_01823_),
    .A2(_02357_),
    .ZN(_02358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08051_ (.I(_01820_),
    .Z(_02359_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08052_ (.A1(_02356_),
    .A2(\mod.u_cpu.rf_ram.memory[70][0] ),
    .B(_02358_),
    .C(_02359_),
    .ZN(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08053_ (.I(_01528_),
    .Z(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08054_ (.A1(_02352_),
    .A2(_02355_),
    .B(_02360_),
    .C(_02361_),
    .ZN(_02362_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08055_ (.I(_01586_),
    .Z(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08056_ (.A1(_02348_),
    .A2(_02351_),
    .B(_02362_),
    .C(_02363_),
    .ZN(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08057_ (.I(_02347_),
    .Z(_02365_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08058_ (.I(_02058_),
    .Z(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08059_ (.I(_01524_),
    .Z(_02367_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08060_ (.I0(\mod.u_cpu.rf_ram.memory[72][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[73][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[74][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[75][0] ),
    .S0(_02366_),
    .S1(_02367_),
    .Z(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08061_ (.I(_01644_),
    .Z(_02369_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08062_ (.I(\mod.u_cpu.rf_ram.memory[77][0] ),
    .ZN(_02370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08063_ (.A1(_02369_),
    .A2(_02370_),
    .ZN(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08064_ (.A1(_02302_),
    .A2(\mod.u_cpu.rf_ram.memory[76][0] ),
    .B(_02371_),
    .ZN(_02372_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08065_ (.I(\mod.u_cpu.rf_ram.memory[79][0] ),
    .ZN(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08066_ (.A1(_01823_),
    .A2(_02373_),
    .ZN(_02374_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08067_ (.A1(_02356_),
    .A2(\mod.u_cpu.rf_ram.memory[78][0] ),
    .B(_02374_),
    .C(_02359_),
    .ZN(_02375_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08068_ (.A1(_02352_),
    .A2(_02372_),
    .B(_02375_),
    .C(_02361_),
    .ZN(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08069_ (.I(_01551_),
    .Z(_02377_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08070_ (.A1(_02365_),
    .A2(_02368_),
    .B(_02376_),
    .C(_02377_),
    .ZN(_02378_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08071_ (.A1(_02149_),
    .A2(_02364_),
    .A3(_02378_),
    .ZN(_02379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08072_ (.I(_01485_),
    .Z(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08073_ (.A1(_02337_),
    .A2(_02346_),
    .B(_02379_),
    .C(_02380_),
    .ZN(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08074_ (.A1(_01483_),
    .A2(_02336_),
    .A3(_02381_),
    .ZN(_02382_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08075_ (.I(_01524_),
    .Z(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08076_ (.I0(\mod.u_cpu.rf_ram.memory[4][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[5][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[6][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[7][0] ),
    .S0(_02366_),
    .S1(_02383_),
    .Z(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08077_ (.I(_01924_),
    .Z(_02385_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08078_ (.I(_01581_),
    .Z(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08079_ (.I0(\mod.u_cpu.rf_ram.memory[0][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[1][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[2][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[3][0] ),
    .S0(_02385_),
    .S1(_02386_),
    .Z(_02387_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08080_ (.I(_02126_),
    .Z(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08081_ (.I0(\mod.u_cpu.rf_ram.memory[12][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[13][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[14][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[15][0] ),
    .S0(_02266_),
    .S1(_02388_),
    .Z(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08082_ (.I0(\mod.u_cpu.rf_ram.memory[8][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[9][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[10][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[11][0] ),
    .S0(_02171_),
    .S1(_02267_),
    .Z(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08083_ (.I(_01679_),
    .Z(_02391_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08084_ (.I0(_02384_),
    .I1(_02387_),
    .I2(_02389_),
    .I3(_02390_),
    .S0(_02391_),
    .S1(_01720_),
    .Z(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08085_ (.I(_02126_),
    .Z(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08086_ (.I0(\mod.u_cpu.rf_ram.memory[24][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[25][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[26][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[27][0] ),
    .S0(_02349_),
    .S1(_02393_),
    .Z(_02394_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08087_ (.I(\mod.u_cpu.rf_ram.memory[29][0] ),
    .ZN(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08088_ (.A1(_02369_),
    .A2(_02395_),
    .ZN(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08089_ (.A1(_02302_),
    .A2(\mod.u_cpu.rf_ram.memory[28][0] ),
    .B(_02396_),
    .ZN(_02397_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08090_ (.I(\mod.u_cpu.rf_ram.memory[31][0] ),
    .ZN(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08091_ (.A1(_01823_),
    .A2(_02398_),
    .ZN(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08092_ (.A1(_02356_),
    .A2(\mod.u_cpu.rf_ram.memory[30][0] ),
    .B(_02399_),
    .C(_02359_),
    .ZN(_02400_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08093_ (.A1(_02352_),
    .A2(_02397_),
    .B(_02400_),
    .C(_02361_),
    .ZN(_02401_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08094_ (.A1(_02348_),
    .A2(_02394_),
    .B(_02401_),
    .C(_02185_),
    .ZN(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08095_ (.I(_01856_),
    .Z(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08096_ (.I0(\mod.u_cpu.rf_ram.memory[16][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[17][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[18][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[19][0] ),
    .S0(_02403_),
    .S1(_02367_),
    .Z(_02404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08097_ (.I(_02154_),
    .Z(_02405_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08098_ (.I(_01644_),
    .Z(_02406_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08099_ (.I(\mod.u_cpu.rf_ram.memory[21][0] ),
    .ZN(_02407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08100_ (.A1(_02406_),
    .A2(_02407_),
    .ZN(_02408_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08101_ (.A1(_02316_),
    .A2(\mod.u_cpu.rf_ram.memory[20][0] ),
    .B(_02408_),
    .ZN(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08102_ (.I(_01646_),
    .Z(_02410_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08103_ (.I(_01778_),
    .Z(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08104_ (.I(\mod.u_cpu.rf_ram.memory[23][0] ),
    .ZN(_02412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08105_ (.A1(_02411_),
    .A2(_02412_),
    .ZN(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08106_ (.A1(_02410_),
    .A2(\mod.u_cpu.rf_ram.memory[22][0] ),
    .B(_02413_),
    .C(_01830_),
    .ZN(_02414_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08107_ (.I(_01765_),
    .Z(_02415_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08108_ (.A1(_02405_),
    .A2(_02409_),
    .B(_02414_),
    .C(_02415_),
    .ZN(_02416_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08109_ (.A1(_02150_),
    .A2(_02404_),
    .B(_02416_),
    .C(_02363_),
    .ZN(_02417_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08110_ (.A1(_01592_),
    .A2(_02402_),
    .A3(_02417_),
    .ZN(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08111_ (.A1(_01693_),
    .A2(_02392_),
    .B(_02418_),
    .C(_02380_),
    .ZN(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08112_ (.I0(\mod.u_cpu.rf_ram.memory[52][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[53][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[54][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[55][0] ),
    .S0(_02403_),
    .S1(_02152_),
    .Z(_02420_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08113_ (.I(_01919_),
    .Z(_02421_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08114_ (.I0(\mod.u_cpu.rf_ram.memory[48][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[49][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[50][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[51][0] ),
    .S0(_02421_),
    .S1(_02350_),
    .Z(_02422_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08115_ (.I0(\mod.u_cpu.rf_ram.memory[60][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[61][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[62][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[63][0] ),
    .S0(_02369_),
    .S1(_02218_),
    .Z(_02423_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08116_ (.I0(\mod.u_cpu.rf_ram.memory[56][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[57][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[58][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[59][0] ),
    .S0(_02242_),
    .S1(_02267_),
    .Z(_02424_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08117_ (.I0(_02420_),
    .I1(_02422_),
    .I2(_02423_),
    .I3(_02424_),
    .S0(_02391_),
    .S1(_01552_),
    .Z(_02425_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08118_ (.I0(\mod.u_cpu.rf_ram.memory[32][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[33][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[34][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[35][0] ),
    .S0(_02403_),
    .S1(_02383_),
    .Z(_02426_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08119_ (.I(\mod.u_cpu.rf_ram.memory[37][0] ),
    .ZN(_02427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08120_ (.A1(_02406_),
    .A2(_02427_),
    .ZN(_02428_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08121_ (.A1(_02329_),
    .A2(\mod.u_cpu.rf_ram.memory[36][0] ),
    .B(_02428_),
    .ZN(_02429_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08122_ (.I(\mod.u_cpu.rf_ram.memory[39][0] ),
    .ZN(_02430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08123_ (.A1(_02411_),
    .A2(_02430_),
    .ZN(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08124_ (.A1(_02410_),
    .A2(\mod.u_cpu.rf_ram.memory[38][0] ),
    .B(_02431_),
    .C(_01828_),
    .ZN(_02432_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08125_ (.A1(_02405_),
    .A2(_02429_),
    .B(_02432_),
    .C(_02415_),
    .ZN(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08126_ (.A1(_02365_),
    .A2(_02426_),
    .B(_02433_),
    .C(_02168_),
    .ZN(_02434_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08127_ (.I0(\mod.u_cpu.rf_ram.memory[40][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[41][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[42][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[43][0] ),
    .S0(_02151_),
    .S1(_02383_),
    .Z(_02435_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08128_ (.I(\mod.u_cpu.rf_ram.memory[45][0] ),
    .ZN(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08129_ (.A1(_02157_),
    .A2(_02436_),
    .ZN(_02437_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08130_ (.A1(_02156_),
    .A2(\mod.u_cpu.rf_ram.memory[44][0] ),
    .B(_02437_),
    .ZN(_02438_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08131_ (.I(\mod.u_cpu.rf_ram.memory[47][0] ),
    .ZN(_02439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08132_ (.A1(_01819_),
    .A2(_02439_),
    .ZN(_02440_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08133_ (.A1(_02161_),
    .A2(\mod.u_cpu.rf_ram.memory[46][0] ),
    .B(_02440_),
    .C(_01828_),
    .ZN(_02441_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08134_ (.A1(_02155_),
    .A2(_02438_),
    .B(_02441_),
    .C(_02166_),
    .ZN(_02442_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08135_ (.A1(_02150_),
    .A2(_02435_),
    .B(_02442_),
    .C(_02185_),
    .ZN(_02443_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08136_ (.A1(_02149_),
    .A2(_02434_),
    .A3(_02443_),
    .ZN(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08137_ (.A1(_02337_),
    .A2(_02425_),
    .B(_02444_),
    .C(_01591_),
    .ZN(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08138_ (.A1(_01475_),
    .A2(_02419_),
    .A3(_02445_),
    .ZN(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08139_ (.A1(_01471_),
    .A2(_02382_),
    .A3(_02446_),
    .ZN(_02447_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08140_ (.A1(_01469_),
    .A2(_02281_),
    .A3(_02447_),
    .Z(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08141_ (.I(_02124_),
    .Z(_02449_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08142_ (.I(_02209_),
    .Z(_02450_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08143_ (.I(_02152_),
    .Z(_02451_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08144_ (.I0(\mod.u_cpu.rf_ram.memory[544][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[545][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[546][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[547][0] ),
    .S0(_02450_),
    .S1(_02451_),
    .Z(_02452_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08145_ (.I(_01782_),
    .Z(_02453_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08146_ (.I(_02453_),
    .Z(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08147_ (.I(_02454_),
    .Z(_02455_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08148_ (.I(_02129_),
    .Z(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08149_ (.I(_01634_),
    .Z(_02457_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08150_ (.I(\mod.u_cpu.rf_ram.memory[549][0] ),
    .ZN(_02458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08151_ (.A1(_02457_),
    .A2(_02458_),
    .ZN(_02459_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08152_ (.A1(_02456_),
    .A2(\mod.u_cpu.rf_ram.memory[548][0] ),
    .B(_02459_),
    .ZN(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08153_ (.I(_02115_),
    .Z(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08154_ (.I(_02116_),
    .Z(_02462_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08155_ (.I(\mod.u_cpu.rf_ram.memory[551][0] ),
    .ZN(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08156_ (.A1(_02462_),
    .A2(_02463_),
    .ZN(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08157_ (.I(_01747_),
    .Z(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08158_ (.A1(_02461_),
    .A2(\mod.u_cpu.rf_ram.memory[550][0] ),
    .B(_02464_),
    .C(_02465_),
    .ZN(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08159_ (.I(_02120_),
    .Z(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08160_ (.A1(_02455_),
    .A2(_02460_),
    .B(_02466_),
    .C(_02467_),
    .ZN(_02468_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08161_ (.I(_02143_),
    .Z(_02469_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08162_ (.A1(_02449_),
    .A2(_02452_),
    .B(_02468_),
    .C(_02469_),
    .ZN(_02470_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08163_ (.I(_01688_),
    .Z(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08164_ (.I(_02329_),
    .Z(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08165_ (.I(_02388_),
    .Z(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08166_ (.I0(\mod.u_cpu.rf_ram.memory[552][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[553][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[554][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[555][0] ),
    .S0(_02472_),
    .S1(_02473_),
    .Z(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08167_ (.I(_01702_),
    .Z(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08168_ (.I(_02475_),
    .Z(_02476_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08169_ (.I(_02047_),
    .Z(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08170_ (.I(_02477_),
    .Z(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08171_ (.I(_01925_),
    .Z(_02479_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08172_ (.I(\mod.u_cpu.rf_ram.memory[557][0] ),
    .ZN(_02480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08173_ (.A1(_02479_),
    .A2(_02480_),
    .ZN(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08174_ (.A1(_02478_),
    .A2(\mod.u_cpu.rf_ram.memory[556][0] ),
    .B(_02481_),
    .ZN(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08175_ (.I(_02175_),
    .Z(_02483_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08176_ (.I(_01745_),
    .Z(_02484_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08177_ (.I(\mod.u_cpu.rf_ram.memory[559][0] ),
    .ZN(_02485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08178_ (.A1(_02484_),
    .A2(_02485_),
    .ZN(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08179_ (.I(_02010_),
    .Z(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08180_ (.A1(_02483_),
    .A2(\mod.u_cpu.rf_ram.memory[558][0] ),
    .B(_02486_),
    .C(_02487_),
    .ZN(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08181_ (.I(_01717_),
    .Z(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08182_ (.A1(_02476_),
    .A2(_02482_),
    .B(_02488_),
    .C(_02489_),
    .ZN(_02490_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08183_ (.I(_02321_),
    .Z(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08184_ (.A1(_02471_),
    .A2(_02474_),
    .B(_02490_),
    .C(_02491_),
    .ZN(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08185_ (.A1(_02470_),
    .A2(_02492_),
    .B(_01447_),
    .ZN(_02493_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08186_ (.I(_01705_),
    .Z(_02494_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08187_ (.I(_02393_),
    .Z(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08188_ (.I0(\mod.u_cpu.rf_ram.memory[568][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[569][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[570][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[571][0] ),
    .S0(_02494_),
    .S1(_02495_),
    .Z(_02496_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08189_ (.I(\mod.u_cpu.rf_ram.memory[573][0] ),
    .ZN(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08190_ (.A1(_02457_),
    .A2(_02497_),
    .ZN(_02498_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08191_ (.A1(_02456_),
    .A2(\mod.u_cpu.rf_ram.memory[572][0] ),
    .B(_02498_),
    .ZN(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08192_ (.I(_02216_),
    .Z(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08193_ (.I(\mod.u_cpu.rf_ram.memory[575][0] ),
    .ZN(_02501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08194_ (.A1(_02500_),
    .A2(_02501_),
    .ZN(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08195_ (.A1(_02461_),
    .A2(\mod.u_cpu.rf_ram.memory[574][0] ),
    .B(_02502_),
    .C(_02465_),
    .ZN(_02503_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08196_ (.A1(_02455_),
    .A2(_02499_),
    .B(_02503_),
    .C(_02467_),
    .ZN(_02504_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08197_ (.I(_02122_),
    .Z(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08198_ (.A1(_02449_),
    .A2(_02496_),
    .B(_02504_),
    .C(_02505_),
    .ZN(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08199_ (.I(_02209_),
    .Z(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08200_ (.I0(\mod.u_cpu.rf_ram.memory[560][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[561][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[562][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[563][0] ),
    .S0(_02507_),
    .S1(_02473_),
    .Z(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08201_ (.I(_01682_),
    .Z(_02509_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08202_ (.I(\mod.u_cpu.rf_ram.memory[565][0] ),
    .ZN(_02510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08203_ (.A1(_02509_),
    .A2(_02510_),
    .ZN(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08204_ (.A1(_02478_),
    .A2(\mod.u_cpu.rf_ram.memory[564][0] ),
    .B(_02511_),
    .ZN(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08205_ (.I(\mod.u_cpu.rf_ram.memory[567][0] ),
    .ZN(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08206_ (.A1(_02484_),
    .A2(_02513_),
    .ZN(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08207_ (.I(_02306_),
    .Z(_02515_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08208_ (.A1(_02483_),
    .A2(\mod.u_cpu.rf_ram.memory[566][0] ),
    .B(_02514_),
    .C(_02515_),
    .ZN(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08209_ (.A1(_02476_),
    .A2(_02512_),
    .B(_02516_),
    .C(_02489_),
    .ZN(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08210_ (.I(_02291_),
    .Z(_02518_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08211_ (.A1(_02471_),
    .A2(_02508_),
    .B(_02517_),
    .C(_02518_),
    .ZN(_02519_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08212_ (.I(_01489_),
    .Z(_02520_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08213_ (.A1(_02506_),
    .A2(_02519_),
    .B(_02520_),
    .ZN(_02521_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08214_ (.A1(_02039_),
    .A2(_02493_),
    .A3(_02521_),
    .ZN(_02522_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08215_ (.I(_02097_),
    .Z(_02523_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08216_ (.I0(\mod.u_cpu.rf_ram.memory[512][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[513][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[514][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[515][0] ),
    .S0(_02494_),
    .S1(_02495_),
    .Z(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08217_ (.I(_02454_),
    .Z(_02525_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08218_ (.I(_02084_),
    .Z(_02526_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08219_ (.I(_02526_),
    .Z(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08220_ (.I(_01538_),
    .Z(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08221_ (.I(\mod.u_cpu.rf_ram.memory[517][0] ),
    .ZN(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08222_ (.A1(_02528_),
    .A2(_02529_),
    .ZN(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08223_ (.A1(_02527_),
    .A2(\mod.u_cpu.rf_ram.memory[516][0] ),
    .B(_02530_),
    .ZN(_02531_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08224_ (.I(_01635_),
    .Z(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08225_ (.I(_02532_),
    .Z(_02533_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08226_ (.I(_02216_),
    .Z(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08227_ (.I(\mod.u_cpu.rf_ram.memory[519][0] ),
    .ZN(_02535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08228_ (.A1(_02534_),
    .A2(_02535_),
    .ZN(_02536_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08229_ (.I(_01747_),
    .Z(_02537_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08230_ (.A1(_02533_),
    .A2(\mod.u_cpu.rf_ram.memory[518][0] ),
    .B(_02536_),
    .C(_02537_),
    .ZN(_02538_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08231_ (.I(_02120_),
    .Z(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08232_ (.A1(_02525_),
    .A2(_02531_),
    .B(_02538_),
    .C(_02539_),
    .ZN(_02540_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08233_ (.A1(_02523_),
    .A2(_02524_),
    .B(_02540_),
    .C(_02469_),
    .ZN(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08234_ (.I(_01688_),
    .Z(_02542_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08235_ (.I(_01855_),
    .Z(_02543_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08236_ (.I0(\mod.u_cpu.rf_ram.memory[520][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[521][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[522][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[523][0] ),
    .S0(_02507_),
    .S1(_02543_),
    .Z(_02544_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08237_ (.I(_02325_),
    .Z(_02545_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08238_ (.I(_02477_),
    .Z(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08239_ (.I(\mod.u_cpu.rf_ram.memory[525][0] ),
    .ZN(_02547_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08240_ (.A1(_02509_),
    .A2(_02547_),
    .ZN(_02548_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08241_ (.A1(_02546_),
    .A2(\mod.u_cpu.rf_ram.memory[524][0] ),
    .B(_02548_),
    .ZN(_02549_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08242_ (.I(_02156_),
    .Z(_02550_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08243_ (.I(_01863_),
    .Z(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08244_ (.I(\mod.u_cpu.rf_ram.memory[527][0] ),
    .ZN(_02552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08245_ (.A1(_02551_),
    .A2(_02552_),
    .ZN(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08246_ (.A1(_02550_),
    .A2(\mod.u_cpu.rf_ram.memory[526][0] ),
    .B(_02553_),
    .C(_02515_),
    .ZN(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08247_ (.I(_02308_),
    .Z(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08248_ (.A1(_02545_),
    .A2(_02549_),
    .B(_02554_),
    .C(_02555_),
    .ZN(_02556_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08249_ (.A1(_02542_),
    .A2(_02544_),
    .B(_02556_),
    .C(_02491_),
    .ZN(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08250_ (.A1(_02541_),
    .A2(_02557_),
    .B(_01447_),
    .ZN(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08251_ (.I(_01757_),
    .Z(_02559_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08252_ (.I(_02559_),
    .Z(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08253_ (.I(_02107_),
    .Z(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08254_ (.I0(\mod.u_cpu.rf_ram.memory[528][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[529][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[530][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[531][0] ),
    .S0(_02560_),
    .S1(_02561_),
    .Z(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08255_ (.I(\mod.u_cpu.rf_ram.memory[533][0] ),
    .ZN(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08256_ (.A1(_02528_),
    .A2(_02563_),
    .ZN(_02564_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08257_ (.A1(_02527_),
    .A2(\mod.u_cpu.rf_ram.memory[532][0] ),
    .B(_02564_),
    .ZN(_02565_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08258_ (.I(_02245_),
    .Z(_02566_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08259_ (.I(\mod.u_cpu.rf_ram.memory[535][0] ),
    .ZN(_02567_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08260_ (.A1(_02566_),
    .A2(_02567_),
    .ZN(_02568_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08261_ (.A1(_02533_),
    .A2(\mod.u_cpu.rf_ram.memory[534][0] ),
    .B(_02568_),
    .C(_02537_),
    .ZN(_02569_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08262_ (.A1(_02525_),
    .A2(_02565_),
    .B(_02569_),
    .C(_02539_),
    .ZN(_02570_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08263_ (.A1(_02523_),
    .A2(_02562_),
    .B(_02570_),
    .C(_02469_),
    .ZN(_02571_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08264_ (.I0(\mod.u_cpu.rf_ram.memory[536][0] ),
    .I1(\mod.u_cpu.rf_ram.memory[537][0] ),
    .I2(\mod.u_cpu.rf_ram.memory[538][0] ),
    .I3(\mod.u_cpu.rf_ram.memory[539][0] ),
    .S0(_02450_),
    .S1(_02451_),
    .Z(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08265_ (.I(\mod.u_cpu.rf_ram.memory[541][0] ),
    .ZN(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08266_ (.A1(_02472_),
    .A2(_02573_),
    .ZN(_02574_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08267_ (.A1(_02546_),
    .A2(\mod.u_cpu.rf_ram.memory[540][0] ),
    .B(_02574_),
    .ZN(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08268_ (.I(\mod.u_cpu.rf_ram.memory[543][0] ),
    .ZN(_02576_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08269_ (.A1(_02551_),
    .A2(_02576_),
    .ZN(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08270_ (.I(_02139_),
    .Z(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08271_ (.A1(_02550_),
    .A2(\mod.u_cpu.rf_ram.memory[542][0] ),
    .B(_02577_),
    .C(_02578_),
    .ZN(_02579_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08272_ (.A1(_02545_),
    .A2(_02575_),
    .B(_02579_),
    .C(_02555_),
    .ZN(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08273_ (.A1(_02542_),
    .A2(_02572_),
    .B(_02580_),
    .C(_02491_),
    .ZN(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08274_ (.A1(_02571_),
    .A2(_02581_),
    .B(_02520_),
    .ZN(_02582_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08275_ (.A1(_01459_),
    .A2(_02558_),
    .A3(_02582_),
    .ZN(_02583_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _08276_ (.A1(_01464_),
    .A2(_01465_),
    .A3(_02522_),
    .A4(_02583_),
    .Z(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _08277_ (.A1(_01466_),
    .A2(_02038_),
    .A3(_02448_),
    .B(_02584_),
    .ZN(_00000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08278_ (.I(_01636_),
    .Z(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08279_ (.I0(\mod.u_cpu.rf_ram.memory[462][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[463][1] ),
    .S(_02585_),
    .Z(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08280_ (.I(\mod.u_cpu.rf_ram.memory[461][1] ),
    .ZN(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08281_ (.A1(_02198_),
    .A2(\mod.u_cpu.rf_ram.memory[460][1] ),
    .ZN(_02588_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08282_ (.A1(_02560_),
    .A2(_02587_),
    .B(_02588_),
    .C(_02188_),
    .ZN(_02589_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08283_ (.A1(_02561_),
    .A2(_02586_),
    .B(_02589_),
    .C(_02080_),
    .ZN(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08284_ (.I(_01851_),
    .Z(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08285_ (.I(_02591_),
    .Z(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08286_ (.I(_02116_),
    .Z(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08287_ (.I(_02030_),
    .Z(_02594_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08288_ (.I0(\mod.u_cpu.rf_ram.memory[456][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[457][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[458][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[459][1] ),
    .S0(_02593_),
    .S1(_02594_),
    .Z(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08289_ (.A1(_02592_),
    .A2(_02595_),
    .B(_02077_),
    .ZN(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08290_ (.I(_01882_),
    .Z(_02597_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08291_ (.I0(\mod.u_cpu.rf_ram.memory[448][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[449][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[450][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[451][1] ),
    .S0(_01508_),
    .S1(_02597_),
    .Z(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08292_ (.I(\mod.u_cpu.rf_ram.memory[453][1] ),
    .ZN(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08293_ (.A1(_01607_),
    .A2(_02599_),
    .ZN(_02600_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08294_ (.A1(_02585_),
    .A2(\mod.u_cpu.rf_ram.memory[452][1] ),
    .B(_02600_),
    .ZN(_02601_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08295_ (.I(\mod.u_cpu.rf_ram.memory[455][1] ),
    .ZN(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08296_ (.A1(_02066_),
    .A2(_02602_),
    .ZN(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08297_ (.A1(_02191_),
    .A2(\mod.u_cpu.rf_ram.memory[454][1] ),
    .B(_02603_),
    .C(_02093_),
    .ZN(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08298_ (.A1(_02487_),
    .A2(_02601_),
    .B(_02604_),
    .C(_02196_),
    .ZN(_02605_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08299_ (.I(_01533_),
    .Z(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08300_ (.A1(_02083_),
    .A2(_02598_),
    .B(_02605_),
    .C(_02606_),
    .ZN(_02607_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08301_ (.A1(_02590_),
    .A2(_02596_),
    .B(_02102_),
    .C(_02607_),
    .ZN(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08302_ (.I(_02040_),
    .Z(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08303_ (.I0(\mod.u_cpu.rf_ram.memory[472][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[473][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[474][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[475][1] ),
    .S0(_02593_),
    .S1(_02454_),
    .Z(_02610_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08304_ (.I(_02350_),
    .Z(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08305_ (.I(\mod.u_cpu.rf_ram.memory[477][1] ),
    .ZN(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08306_ (.A1(_02593_),
    .A2(_02612_),
    .ZN(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08307_ (.A1(_02566_),
    .A2(\mod.u_cpu.rf_ram.memory[476][1] ),
    .B(_02613_),
    .ZN(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08308_ (.I(\mod.u_cpu.rf_ram.memory[479][1] ),
    .ZN(_02615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08309_ (.A1(_02532_),
    .A2(_02615_),
    .ZN(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08310_ (.A1(_02198_),
    .A2(\mod.u_cpu.rf_ram.memory[478][1] ),
    .B(_02616_),
    .C(_01751_),
    .ZN(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08311_ (.A1(_02611_),
    .A2(_02614_),
    .B(_02617_),
    .C(_01742_),
    .ZN(_02618_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08312_ (.A1(_02592_),
    .A2(_02610_),
    .B(_02618_),
    .C(_01678_),
    .ZN(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08313_ (.I0(\mod.u_cpu.rf_ram.memory[464][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[465][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[466][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[467][1] ),
    .S0(_02593_),
    .S1(_02454_),
    .Z(_02620_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08314_ (.I(\mod.u_cpu.rf_ram.memory[469][1] ),
    .ZN(_02621_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08315_ (.A1(_02225_),
    .A2(_02621_),
    .ZN(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08316_ (.A1(_02566_),
    .A2(\mod.u_cpu.rf_ram.memory[468][1] ),
    .B(_02622_),
    .ZN(_02623_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08317_ (.I(\mod.u_cpu.rf_ram.memory[471][1] ),
    .ZN(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08318_ (.A1(_02115_),
    .A2(_02624_),
    .ZN(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08319_ (.A1(_02198_),
    .A2(\mod.u_cpu.rf_ram.memory[470][1] ),
    .B(_02625_),
    .C(_01751_),
    .ZN(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08320_ (.A1(_02611_),
    .A2(_02623_),
    .B(_02626_),
    .C(_01742_),
    .ZN(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08321_ (.A1(_02592_),
    .A2(_02620_),
    .B(_02627_),
    .C(_01658_),
    .ZN(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08322_ (.A1(_02609_),
    .A2(_02619_),
    .A3(_02628_),
    .ZN(_02629_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08323_ (.A1(_02039_),
    .A2(_02608_),
    .A3(_02629_),
    .ZN(_02630_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08324_ (.I(_02347_),
    .Z(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08325_ (.I(_01495_),
    .Z(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08326_ (.I(_01637_),
    .Z(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08327_ (.I0(\mod.u_cpu.rf_ram.memory[496][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[497][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[498][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[499][1] ),
    .S0(_02632_),
    .S1(_02633_),
    .Z(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08328_ (.I(\mod.u_cpu.rf_ram.memory[501][1] ),
    .ZN(_02635_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08329_ (.A1(_02421_),
    .A2(_02635_),
    .ZN(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08330_ (.A1(_02559_),
    .A2(\mod.u_cpu.rf_ram.memory[500][1] ),
    .B(_02636_),
    .ZN(_02637_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08331_ (.I(_01537_),
    .Z(_02638_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08332_ (.I(\mod.u_cpu.rf_ram.memory[503][1] ),
    .ZN(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08333_ (.A1(_02197_),
    .A2(_02639_),
    .ZN(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08334_ (.A1(_02638_),
    .A2(\mod.u_cpu.rf_ram.memory[502][1] ),
    .B(_02640_),
    .C(_01615_),
    .ZN(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08335_ (.A1(_02597_),
    .A2(_02637_),
    .B(_02641_),
    .C(_01651_),
    .ZN(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08336_ (.A1(_02631_),
    .A2(_02634_),
    .B(_02642_),
    .C(_01587_),
    .ZN(_02643_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08337_ (.I0(\mod.u_cpu.rf_ram.memory[504][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[505][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[506][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[507][1] ),
    .S0(_02385_),
    .S1(_02633_),
    .Z(_02644_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08338_ (.I(\mod.u_cpu.rf_ram.memory[509][1] ),
    .ZN(_02645_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08339_ (.A1(_02421_),
    .A2(_02645_),
    .ZN(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08340_ (.A1(_02559_),
    .A2(\mod.u_cpu.rf_ram.memory[508][1] ),
    .B(_02646_),
    .ZN(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08341_ (.I(\mod.u_cpu.rf_ram.memory[511][1] ),
    .ZN(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08342_ (.A1(_02220_),
    .A2(_02648_),
    .ZN(_02649_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08343_ (.A1(_02638_),
    .A2(\mod.u_cpu.rf_ram.memory[510][1] ),
    .B(_02649_),
    .C(_01821_),
    .ZN(_02650_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08344_ (.A1(_02597_),
    .A2(_02647_),
    .B(_02650_),
    .C(_01651_),
    .ZN(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08345_ (.A1(_02631_),
    .A2(_02644_),
    .B(_02651_),
    .C(_02377_),
    .ZN(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08346_ (.A1(_01592_),
    .A2(_02643_),
    .A3(_02652_),
    .ZN(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08347_ (.I(_02218_),
    .Z(_02654_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08348_ (.I0(\mod.u_cpu.rf_ram.memory[494][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[495][1] ),
    .S(_01709_),
    .Z(_02655_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08349_ (.I(_01841_),
    .Z(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08350_ (.I(\mod.u_cpu.rf_ram.memory[493][1] ),
    .ZN(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08351_ (.A1(_02085_),
    .A2(\mod.u_cpu.rf_ram.memory[492][1] ),
    .ZN(_02658_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08352_ (.A1(_02656_),
    .A2(_02657_),
    .B(_02658_),
    .C(_02067_),
    .ZN(_02659_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08353_ (.I(_01679_),
    .Z(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08354_ (.A1(_02654_),
    .A2(_02655_),
    .B(_02659_),
    .C(_02660_),
    .ZN(_02661_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08355_ (.I0(\mod.u_cpu.rf_ram.memory[488][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[489][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[490][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[491][1] ),
    .S0(_02385_),
    .S1(_02633_),
    .Z(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08356_ (.A1(_02631_),
    .A2(_02662_),
    .B(_01618_),
    .ZN(_02663_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08357_ (.I(_01890_),
    .Z(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08358_ (.I(_01991_),
    .Z(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08359_ (.I(_01762_),
    .Z(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08360_ (.I0(\mod.u_cpu.rf_ram.memory[480][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[481][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[482][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[483][1] ),
    .S0(_01963_),
    .S1(_02666_),
    .Z(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08361_ (.I(_01960_),
    .Z(_02668_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08362_ (.I(\mod.u_cpu.rf_ram.memory[485][1] ),
    .ZN(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08363_ (.A1(_01561_),
    .A2(_02669_),
    .ZN(_02670_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08364_ (.A1(_02638_),
    .A2(\mod.u_cpu.rf_ram.memory[484][1] ),
    .B(_02670_),
    .ZN(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08365_ (.I(_02026_),
    .Z(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08366_ (.I(\mod.u_cpu.rf_ram.memory[487][1] ),
    .ZN(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08367_ (.A1(_02672_),
    .A2(_02673_),
    .ZN(_02674_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08368_ (.A1(_01567_),
    .A2(\mod.u_cpu.rf_ram.memory[486][1] ),
    .B(_02674_),
    .C(_02109_),
    .ZN(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08369_ (.A1(_02668_),
    .A2(_02671_),
    .B(_02675_),
    .C(_01687_),
    .ZN(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08370_ (.I(_01886_),
    .Z(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08371_ (.A1(_02665_),
    .A2(_02667_),
    .B(_02676_),
    .C(_02677_),
    .ZN(_02678_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08372_ (.A1(_02661_),
    .A2(_02663_),
    .B(_02664_),
    .C(_02678_),
    .ZN(_02679_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08373_ (.A1(_01591_),
    .A2(_02653_),
    .A3(_02679_),
    .ZN(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08374_ (.A1(_02148_),
    .A2(_02680_),
    .Z(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08375_ (.I0(\mod.u_cpu.rf_ram.memory[430][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[431][1] ),
    .S(_02585_),
    .Z(_02682_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08376_ (.I(\mod.u_cpu.rf_ram.memory[429][1] ),
    .ZN(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08377_ (.A1(_02656_),
    .A2(\mod.u_cpu.rf_ram.memory[428][1] ),
    .ZN(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08378_ (.A1(_02560_),
    .A2(_02683_),
    .B(_02684_),
    .C(_02594_),
    .ZN(_02685_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08379_ (.A1(_02561_),
    .A2(_02682_),
    .B(_02685_),
    .C(_02080_),
    .ZN(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08380_ (.I(_02591_),
    .Z(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08381_ (.I(_01879_),
    .Z(_02688_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08382_ (.I0(\mod.u_cpu.rf_ram.memory[424][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[425][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[426][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[427][1] ),
    .S0(_02688_),
    .S1(_02475_),
    .Z(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08383_ (.A1(_02687_),
    .A2(_02689_),
    .B(_02077_),
    .ZN(_02690_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08384_ (.I0(\mod.u_cpu.rf_ram.memory[416][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[417][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[418][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[419][1] ),
    .S0(_02559_),
    .S1(_02155_),
    .Z(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08385_ (.I(_02220_),
    .Z(_02692_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08386_ (.I(\mod.u_cpu.rf_ram.memory[421][1] ),
    .ZN(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08387_ (.A1(_02532_),
    .A2(_02693_),
    .ZN(_02694_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08388_ (.A1(_02692_),
    .A2(\mod.u_cpu.rf_ram.memory[420][1] ),
    .B(_02694_),
    .ZN(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08389_ (.I(\mod.u_cpu.rf_ram.memory[423][1] ),
    .ZN(_02696_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08390_ (.A1(_02272_),
    .A2(_02696_),
    .ZN(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08391_ (.A1(_02191_),
    .A2(\mod.u_cpu.rf_ram.memory[422][1] ),
    .B(_02697_),
    .C(_02323_),
    .ZN(_02698_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08392_ (.A1(_02188_),
    .A2(_02695_),
    .B(_02698_),
    .C(_02196_),
    .ZN(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08393_ (.A1(_02083_),
    .A2(_02691_),
    .B(_02699_),
    .C(_02606_),
    .ZN(_02700_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08394_ (.A1(_02686_),
    .A2(_02690_),
    .B(_02105_),
    .C(_02700_),
    .ZN(_02701_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08395_ (.I0(\mod.u_cpu.rf_ram.memory[432][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[433][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[434][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[435][1] ),
    .S0(_02688_),
    .S1(_02475_),
    .Z(_02702_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08396_ (.I(\mod.u_cpu.rf_ram.memory[437][1] ),
    .ZN(_02703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08397_ (.A1(_02111_),
    .A2(_02703_),
    .ZN(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08398_ (.A1(_02500_),
    .A2(\mod.u_cpu.rf_ram.memory[436][1] ),
    .B(_02704_),
    .ZN(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08399_ (.I(\mod.u_cpu.rf_ram.memory[439][1] ),
    .ZN(_02706_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08400_ (.A1(_01709_),
    .A2(_02706_),
    .ZN(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08401_ (.A1(_02692_),
    .A2(\mod.u_cpu.rf_ram.memory[438][1] ),
    .B(_02707_),
    .C(_01981_),
    .ZN(_02708_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08402_ (.A1(_02654_),
    .A2(_02705_),
    .B(_02708_),
    .C(_01979_),
    .ZN(_02709_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08403_ (.A1(_02687_),
    .A2(_02702_),
    .B(_02709_),
    .C(_02606_),
    .ZN(_02710_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08404_ (.I(_01518_),
    .Z(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08405_ (.I0(\mod.u_cpu.rf_ram.memory[440][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[441][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[442][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[443][1] ),
    .S0(_02711_),
    .S1(_01703_),
    .Z(_02712_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08406_ (.I(\mod.u_cpu.rf_ram.memory[445][1] ),
    .ZN(_02713_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08407_ (.A1(_02111_),
    .A2(_02713_),
    .ZN(_02714_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08408_ (.A1(_02462_),
    .A2(\mod.u_cpu.rf_ram.memory[444][1] ),
    .B(_02714_),
    .ZN(_02715_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08409_ (.I(\mod.u_cpu.rf_ram.memory[447][1] ),
    .ZN(_02716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08410_ (.A1(_01709_),
    .A2(_02716_),
    .ZN(_02717_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08411_ (.A1(_02656_),
    .A2(\mod.u_cpu.rf_ram.memory[446][1] ),
    .B(_02717_),
    .C(_01961_),
    .ZN(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08412_ (.A1(_02654_),
    .A2(_02715_),
    .B(_02718_),
    .C(_01992_),
    .ZN(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08413_ (.A1(_02539_),
    .A2(_02712_),
    .B(_02719_),
    .C(_01678_),
    .ZN(_02720_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08414_ (.A1(_02609_),
    .A2(_02710_),
    .A3(_02720_),
    .ZN(_02721_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08415_ (.A1(_01459_),
    .A2(_02701_),
    .A3(_02721_),
    .ZN(_02722_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08416_ (.I0(\mod.u_cpu.rf_ram.memory[408][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[409][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[410][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[411][1] ),
    .S0(_02225_),
    .S1(_02325_),
    .Z(_02723_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08417_ (.I(\mod.u_cpu.rf_ram.memory[413][1] ),
    .ZN(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08418_ (.A1(_02526_),
    .A2(_02724_),
    .ZN(_02725_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08419_ (.A1(_02534_),
    .A2(\mod.u_cpu.rf_ram.memory[412][1] ),
    .B(_02725_),
    .ZN(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08420_ (.I(\mod.u_cpu.rf_ram.memory[415][1] ),
    .ZN(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08421_ (.A1(_02244_),
    .A2(_02727_),
    .ZN(_02728_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08422_ (.A1(_02692_),
    .A2(\mod.u_cpu.rf_ram.memory[414][1] ),
    .B(_02728_),
    .C(_01773_),
    .ZN(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08423_ (.I(_01914_),
    .Z(_02730_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08424_ (.A1(_02611_),
    .A2(_02726_),
    .B(_02729_),
    .C(_02730_),
    .ZN(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08425_ (.A1(_02687_),
    .A2(_02723_),
    .B(_02731_),
    .C(_01678_),
    .ZN(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08426_ (.I0(\mod.u_cpu.rf_ram.memory[400][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[401][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[402][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[403][1] ),
    .S0(_02688_),
    .S1(_02475_),
    .Z(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08427_ (.I(\mod.u_cpu.rf_ram.memory[405][1] ),
    .ZN(_02734_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08428_ (.A1(_02526_),
    .A2(_02734_),
    .ZN(_02735_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08429_ (.A1(_02534_),
    .A2(\mod.u_cpu.rf_ram.memory[404][1] ),
    .B(_02735_),
    .ZN(_02736_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08430_ (.I(\mod.u_cpu.rf_ram.memory[407][1] ),
    .ZN(_02737_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08431_ (.A1(_02244_),
    .A2(_02737_),
    .ZN(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08432_ (.A1(_02692_),
    .A2(\mod.u_cpu.rf_ram.memory[406][1] ),
    .B(_02738_),
    .C(_01918_),
    .ZN(_02739_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08433_ (.A1(_02654_),
    .A2(_02736_),
    .B(_02739_),
    .C(_02730_),
    .ZN(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08434_ (.A1(_02687_),
    .A2(_02733_),
    .B(_02740_),
    .C(_01658_),
    .ZN(_02741_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08435_ (.A1(_02609_),
    .A2(_02732_),
    .A3(_02741_),
    .ZN(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08436_ (.I0(\mod.u_cpu.rf_ram.memory[384][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[385][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[386][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[387][1] ),
    .S0(_01994_),
    .S1(_02010_),
    .Z(_02743_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08437_ (.A1(_01680_),
    .A2(_02743_),
    .ZN(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08438_ (.I0(\mod.u_cpu.rf_ram.memory[388][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[389][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[390][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[391][1] ),
    .S0(_02020_),
    .S1(_01995_),
    .Z(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08439_ (.A1(_01770_),
    .A2(_02745_),
    .ZN(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08440_ (.A1(_02143_),
    .A2(_02744_),
    .A3(_02746_),
    .ZN(_02747_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08441_ (.I(_01762_),
    .Z(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08442_ (.I0(\mod.u_cpu.rf_ram.memory[392][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[393][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[394][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[395][1] ),
    .S0(_02020_),
    .S1(_02748_),
    .Z(_02749_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08443_ (.A1(_01680_),
    .A2(_02749_),
    .ZN(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08444_ (.I(_01919_),
    .Z(_02751_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08445_ (.I0(\mod.u_cpu.rf_ram.memory[396][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[397][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[398][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[399][1] ),
    .S0(_02751_),
    .S1(_02748_),
    .Z(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08446_ (.A1(_02730_),
    .A2(_02752_),
    .ZN(_02753_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08447_ (.A1(_02230_),
    .A2(_02750_),
    .A3(_02753_),
    .ZN(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08448_ (.A1(_02747_),
    .A2(_02754_),
    .ZN(_02755_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08449_ (.A1(_02337_),
    .A2(_02755_),
    .B(_01591_),
    .ZN(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08450_ (.A1(_02742_),
    .A2(_02756_),
    .B(_01483_),
    .ZN(_02757_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08451_ (.A1(_02630_),
    .A2(_02681_),
    .B1(_02722_),
    .B2(_02757_),
    .ZN(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08452_ (.I(_01615_),
    .Z(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08453_ (.I0(\mod.u_cpu.rf_ram.memory[382][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[383][1] ),
    .S(_02125_),
    .Z(_02760_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08454_ (.I(\mod.u_cpu.rf_ram.memory[381][1] ),
    .ZN(_02761_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08455_ (.A1(_01496_),
    .A2(\mod.u_cpu.rf_ram.memory[380][1] ),
    .ZN(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08456_ (.A1(_02711_),
    .A2(_02761_),
    .B(_02762_),
    .C(_01698_),
    .ZN(_02763_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08457_ (.I(_01660_),
    .Z(_02764_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08458_ (.A1(_02759_),
    .A2(_02760_),
    .B(_02763_),
    .C(_02764_),
    .ZN(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08459_ (.I0(\mod.u_cpu.rf_ram.memory[376][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[377][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[378][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[379][1] ),
    .S0(_01957_),
    .S1(_01958_),
    .Z(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08460_ (.A1(_01956_),
    .A2(_02766_),
    .B(_01788_),
    .ZN(_02767_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08461_ (.I0(\mod.u_cpu.rf_ram.memory[368][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[369][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[370][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[371][1] ),
    .S0(_01837_),
    .S1(_01838_),
    .Z(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08462_ (.I(\mod.u_cpu.rf_ram.memory[373][1] ),
    .ZN(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08463_ (.A1(_01858_),
    .A2(_02769_),
    .ZN(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08464_ (.A1(_02059_),
    .A2(\mod.u_cpu.rf_ram.memory[372][1] ),
    .B(_02770_),
    .ZN(_02771_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08465_ (.I(\mod.u_cpu.rf_ram.memory[375][1] ),
    .ZN(_02772_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08466_ (.A1(_01864_),
    .A2(_02772_),
    .ZN(_02773_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08467_ (.A1(_02303_),
    .A2(\mod.u_cpu.rf_ram.memory[374][1] ),
    .B(_02773_),
    .C(_01867_),
    .ZN(_02774_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08468_ (.A1(_01855_),
    .A2(_02771_),
    .B(_02774_),
    .C(_01631_),
    .ZN(_02775_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08469_ (.A1(_01852_),
    .A2(_02768_),
    .B(_02775_),
    .C(_01887_),
    .ZN(_02776_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08470_ (.A1(_02765_),
    .A2(_02767_),
    .B(_02776_),
    .C(_01849_),
    .ZN(_02777_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08471_ (.I(_01991_),
    .Z(_02778_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08472_ (.I0(\mod.u_cpu.rf_ram.memory[360][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[361][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[362][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[363][1] ),
    .S0(_02751_),
    .S1(_02748_),
    .Z(_02779_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08473_ (.I(\mod.u_cpu.rf_ram.memory[365][1] ),
    .ZN(_02780_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08474_ (.A1(_01729_),
    .A2(_02780_),
    .ZN(_02781_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08475_ (.A1(_02022_),
    .A2(\mod.u_cpu.rf_ram.memory[364][1] ),
    .B(_02781_),
    .ZN(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08476_ (.I(\mod.u_cpu.rf_ram.memory[367][1] ),
    .ZN(_02783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08477_ (.A1(_02027_),
    .A2(_02783_),
    .ZN(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08478_ (.A1(_01875_),
    .A2(\mod.u_cpu.rf_ram.memory[366][1] ),
    .B(_02784_),
    .C(_02030_),
    .ZN(_02785_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08479_ (.A1(_01997_),
    .A2(_02782_),
    .B(_02785_),
    .C(_02096_),
    .ZN(_02786_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08480_ (.A1(_02778_),
    .A2(_02779_),
    .B(_02786_),
    .C(_02007_),
    .ZN(_02787_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08481_ (.I0(\mod.u_cpu.rf_ram.memory[352][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[353][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[354][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[355][1] ),
    .S0(_01920_),
    .S1(_02666_),
    .Z(_02788_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08482_ (.I(\mod.u_cpu.rf_ram.memory[357][1] ),
    .ZN(_02789_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08483_ (.A1(_01520_),
    .A2(_02789_),
    .ZN(_02790_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08484_ (.A1(_02041_),
    .A2(\mod.u_cpu.rf_ram.memory[356][1] ),
    .B(_02790_),
    .ZN(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08485_ (.I(\mod.u_cpu.rf_ram.memory[359][1] ),
    .ZN(_02792_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08486_ (.A1(_02672_),
    .A2(_02792_),
    .ZN(_02793_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08487_ (.A1(_01496_),
    .A2(\mod.u_cpu.rf_ram.memory[358][1] ),
    .B(_02793_),
    .C(_02453_),
    .ZN(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08488_ (.A1(_02668_),
    .A2(_02791_),
    .B(_02794_),
    .C(_02096_),
    .ZN(_02795_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08489_ (.A1(_02778_),
    .A2(_02788_),
    .B(_02795_),
    .C(_02677_),
    .ZN(_02796_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08490_ (.A1(_02664_),
    .A2(_02787_),
    .A3(_02796_),
    .ZN(_02797_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08491_ (.A1(_01848_),
    .A2(_02777_),
    .A3(_02797_),
    .ZN(_02798_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08492_ (.I0(\mod.u_cpu.rf_ram.memory[328][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[329][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[330][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[331][1] ),
    .S0(_01920_),
    .S1(_02666_),
    .Z(_02799_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08493_ (.I(\mod.u_cpu.rf_ram.memory[333][1] ),
    .ZN(_02800_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08494_ (.A1(_01729_),
    .A2(_02800_),
    .ZN(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08495_ (.A1(_02041_),
    .A2(\mod.u_cpu.rf_ram.memory[332][1] ),
    .B(_02801_),
    .ZN(_02802_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08496_ (.I(\mod.u_cpu.rf_ram.memory[335][1] ),
    .ZN(_02803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08497_ (.A1(_02672_),
    .A2(_02803_),
    .ZN(_02804_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08498_ (.A1(_01875_),
    .A2(\mod.u_cpu.rf_ram.memory[334][1] ),
    .B(_02804_),
    .C(_02453_),
    .ZN(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08499_ (.A1(_02668_),
    .A2(_02802_),
    .B(_02805_),
    .C(_02096_),
    .ZN(_02806_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08500_ (.A1(_02778_),
    .A2(_02799_),
    .B(_02806_),
    .C(_01870_),
    .ZN(_02807_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08501_ (.I0(\mod.u_cpu.rf_ram.memory[320][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[321][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[322][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[323][1] ),
    .S0(_01920_),
    .S1(_02666_),
    .Z(_02808_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08502_ (.I(\mod.u_cpu.rf_ram.memory[325][1] ),
    .ZN(_02809_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08503_ (.A1(_01520_),
    .A2(_02809_),
    .ZN(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08504_ (.A1(_02041_),
    .A2(\mod.u_cpu.rf_ram.memory[324][1] ),
    .B(_02810_),
    .ZN(_02811_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08505_ (.I(\mod.u_cpu.rf_ram.memory[327][1] ),
    .ZN(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08506_ (.A1(_02672_),
    .A2(_02812_),
    .ZN(_02813_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08507_ (.A1(_01540_),
    .A2(\mod.u_cpu.rf_ram.memory[326][1] ),
    .B(_02813_),
    .C(_02453_),
    .ZN(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08508_ (.A1(_02668_),
    .A2(_02811_),
    .B(_02814_),
    .C(_01687_),
    .ZN(_02815_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08509_ (.A1(_02665_),
    .A2(_02808_),
    .B(_02815_),
    .C(_02677_),
    .ZN(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08510_ (.A1(_02664_),
    .A2(_02807_),
    .A3(_02816_),
    .ZN(_02817_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08511_ (.I0(\mod.u_cpu.rf_ram.memory[350][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[351][1] ),
    .S(_01664_),
    .Z(_02818_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08512_ (.I(\mod.u_cpu.rf_ram.memory[349][1] ),
    .ZN(_02819_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08513_ (.A1(_01605_),
    .A2(\mod.u_cpu.rf_ram.memory[348][1] ),
    .ZN(_02820_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08514_ (.A1(_02526_),
    .A2(_02819_),
    .B(_02820_),
    .C(_01501_),
    .ZN(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08515_ (.A1(_02759_),
    .A2(_02818_),
    .B(_02821_),
    .C(_02764_),
    .ZN(_02822_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08516_ (.I0(\mod.u_cpu.rf_ram.memory[344][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[345][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[346][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[347][1] ),
    .S0(_02751_),
    .S1(_02748_),
    .Z(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08517_ (.A1(_02778_),
    .A2(_02823_),
    .B(_01788_),
    .ZN(_02824_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08518_ (.I0(\mod.u_cpu.rf_ram.memory[336][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[337][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[338][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[339][1] ),
    .S0(_01841_),
    .S1(_01844_),
    .Z(_02825_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08519_ (.I(\mod.u_cpu.rf_ram.memory[341][1] ),
    .ZN(_02826_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08520_ (.A1(_01858_),
    .A2(_02826_),
    .ZN(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08521_ (.A1(_01893_),
    .A2(\mod.u_cpu.rf_ram.memory[340][1] ),
    .B(_02827_),
    .ZN(_02828_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08522_ (.I(\mod.u_cpu.rf_ram.memory[343][1] ),
    .ZN(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08523_ (.A1(_01864_),
    .A2(_02829_),
    .ZN(_02830_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08524_ (.A1(_01879_),
    .A2(\mod.u_cpu.rf_ram.memory[342][1] ),
    .B(_02830_),
    .C(_01867_),
    .ZN(_02831_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08525_ (.A1(_01874_),
    .A2(_02828_),
    .B(_02831_),
    .C(_01884_),
    .ZN(_02832_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08526_ (.A1(_01872_),
    .A2(_02825_),
    .B(_02832_),
    .C(_01887_),
    .ZN(_02833_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08527_ (.A1(_02822_),
    .A2(_02824_),
    .B(_02040_),
    .C(_02833_),
    .ZN(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08528_ (.A1(_01977_),
    .A2(_02817_),
    .A3(_02834_),
    .ZN(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08529_ (.A1(_02148_),
    .A2(_02798_),
    .A3(_02835_),
    .ZN(_02836_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08530_ (.I0(\mod.u_cpu.rf_ram.memory[302][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[303][1] ),
    .S(_02272_),
    .Z(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08531_ (.I(\mod.u_cpu.rf_ram.memory[301][1] ),
    .ZN(_02838_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08532_ (.A1(_02059_),
    .A2(\mod.u_cpu.rf_ram.memory[300][1] ),
    .ZN(_02839_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08533_ (.A1(_02225_),
    .A2(_02838_),
    .B(_02839_),
    .C(_01683_),
    .ZN(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08534_ (.A1(_02188_),
    .A2(_02837_),
    .B(_02840_),
    .C(_01833_),
    .ZN(_02841_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08535_ (.I0(\mod.u_cpu.rf_ram.memory[296][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[297][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[298][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[299][1] ),
    .S0(_01753_),
    .S1(_01916_),
    .Z(_02842_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08536_ (.A1(_02730_),
    .A2(_02842_),
    .B(_02207_),
    .ZN(_02843_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08537_ (.I0(\mod.u_cpu.rf_ram.memory[288][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[289][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[290][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[291][1] ),
    .S0(_01826_),
    .S1(_02164_),
    .Z(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08538_ (.I(\mod.u_cpu.rf_ram.memory[293][1] ),
    .ZN(_02845_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08539_ (.A1(_01843_),
    .A2(_02845_),
    .ZN(_02846_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08540_ (.A1(_01807_),
    .A2(\mod.u_cpu.rf_ram.memory[292][1] ),
    .B(_02846_),
    .ZN(_02847_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08541_ (.I(\mod.u_cpu.rf_ram.memory[295][1] ),
    .ZN(_02848_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08542_ (.A1(_02091_),
    .A2(_02848_),
    .ZN(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08543_ (.A1(_02216_),
    .A2(\mod.u_cpu.rf_ram.memory[294][1] ),
    .B(_02849_),
    .C(_01504_),
    .ZN(_02850_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08544_ (.A1(_02295_),
    .A2(_02847_),
    .B(_02850_),
    .C(_01492_),
    .ZN(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08545_ (.I(_01886_),
    .Z(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08546_ (.A1(_02196_),
    .A2(_02844_),
    .B(_02851_),
    .C(_02852_),
    .ZN(_02853_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08547_ (.A1(_02841_),
    .A2(_02843_),
    .B(_01891_),
    .C(_02853_),
    .ZN(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08548_ (.I0(\mod.u_cpu.rf_ram.memory[312][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[313][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[314][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[315][1] ),
    .S0(_01802_),
    .S1(_01932_),
    .Z(_02855_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08549_ (.I(\mod.u_cpu.rf_ram.memory[317][1] ),
    .ZN(_02856_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08550_ (.A1(_01934_),
    .A2(_02856_),
    .ZN(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08551_ (.A1(_01962_),
    .A2(\mod.u_cpu.rf_ram.memory[316][1] ),
    .B(_02857_),
    .ZN(_02858_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08552_ (.I(\mod.u_cpu.rf_ram.memory[319][1] ),
    .ZN(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08553_ (.A1(_01949_),
    .A2(_02859_),
    .ZN(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08554_ (.A1(_01938_),
    .A2(\mod.u_cpu.rf_ram.memory[318][1] ),
    .B(_02860_),
    .C(_01952_),
    .ZN(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08555_ (.A1(_01981_),
    .A2(_02858_),
    .B(_02861_),
    .C(_01929_),
    .ZN(_02862_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08556_ (.A1(_01915_),
    .A2(_02855_),
    .B(_02862_),
    .C(_01812_),
    .ZN(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08557_ (.I0(\mod.u_cpu.rf_ram.memory[304][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[305][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[306][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[307][1] ),
    .S0(_01994_),
    .S1(_02010_),
    .Z(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08558_ (.I(\mod.u_cpu.rf_ram.memory[309][1] ),
    .ZN(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08559_ (.A1(_01963_),
    .A2(_02865_),
    .ZN(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08560_ (.A1(_01998_),
    .A2(\mod.u_cpu.rf_ram.memory[308][1] ),
    .B(_02866_),
    .ZN(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08561_ (.I(\mod.u_cpu.rf_ram.memory[311][1] ),
    .ZN(_02868_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08562_ (.A1(_01967_),
    .A2(_02868_),
    .ZN(_02869_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08563_ (.A1(_01697_),
    .A2(\mod.u_cpu.rf_ram.memory[310][1] ),
    .B(_02869_),
    .C(_01970_),
    .ZN(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08564_ (.A1(_01961_),
    .A2(_02867_),
    .B(_02870_),
    .C(_01972_),
    .ZN(_02871_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08565_ (.A1(_01956_),
    .A2(_02864_),
    .B(_02871_),
    .C(_01989_),
    .ZN(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08566_ (.A1(_01791_),
    .A2(_02863_),
    .A3(_02872_),
    .ZN(_02873_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08567_ (.A1(_01848_),
    .A2(_02854_),
    .A3(_02873_),
    .ZN(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08568_ (.I0(\mod.u_cpu.rf_ram.memory[272][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[273][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[274][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[275][1] ),
    .S0(_01957_),
    .S1(_01958_),
    .Z(_02875_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08569_ (.I(\mod.u_cpu.rf_ram.memory[277][1] ),
    .ZN(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08570_ (.A1(_01963_),
    .A2(_02876_),
    .ZN(_02877_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08571_ (.A1(_01962_),
    .A2(\mod.u_cpu.rf_ram.memory[276][1] ),
    .B(_02877_),
    .ZN(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08572_ (.I(\mod.u_cpu.rf_ram.memory[279][1] ),
    .ZN(_02879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08573_ (.A1(_01949_),
    .A2(_02879_),
    .ZN(_02880_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08574_ (.A1(_01697_),
    .A2(\mod.u_cpu.rf_ram.memory[278][1] ),
    .B(_02880_),
    .C(_01952_),
    .ZN(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08575_ (.A1(_01981_),
    .A2(_02878_),
    .B(_02881_),
    .C(_01972_),
    .ZN(_02882_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08576_ (.A1(_01979_),
    .A2(_02875_),
    .B(_02882_),
    .C(_01989_),
    .ZN(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08577_ (.I0(\mod.u_cpu.rf_ram.memory[280][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[281][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[282][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[283][1] ),
    .S0(_02020_),
    .S1(_01995_),
    .Z(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08578_ (.I(\mod.u_cpu.rf_ram.memory[285][1] ),
    .ZN(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08579_ (.A1(_01711_),
    .A2(_02885_),
    .ZN(_02886_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08580_ (.A1(_01998_),
    .A2(\mod.u_cpu.rf_ram.memory[284][1] ),
    .B(_02886_),
    .ZN(_02887_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08581_ (.I(\mod.u_cpu.rf_ram.memory[287][1] ),
    .ZN(_02888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08582_ (.A1(_02027_),
    .A2(_02888_),
    .ZN(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08583_ (.A1(_01722_),
    .A2(\mod.u_cpu.rf_ram.memory[286][1] ),
    .B(_02889_),
    .C(_02030_),
    .ZN(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08584_ (.A1(_01997_),
    .A2(_02887_),
    .B(_02890_),
    .C(_02005_),
    .ZN(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08585_ (.A1(_01992_),
    .A2(_02884_),
    .B(_02891_),
    .C(_02007_),
    .ZN(_02892_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08586_ (.A1(_01978_),
    .A2(_02883_),
    .A3(_02892_),
    .ZN(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08587_ (.I0(\mod.u_cpu.rf_ram.memory[270][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[271][1] ),
    .S(_02106_),
    .Z(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08588_ (.I(\mod.u_cpu.rf_ram.memory[269][1] ),
    .ZN(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08589_ (.A1(_01496_),
    .A2(\mod.u_cpu.rf_ram.memory[268][1] ),
    .ZN(_02896_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08590_ (.A1(_02688_),
    .A2(_02895_),
    .B(_02896_),
    .C(_01698_),
    .ZN(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08591_ (.A1(_02759_),
    .A2(_02894_),
    .B(_02897_),
    .C(_02764_),
    .ZN(_02898_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08592_ (.I0(\mod.u_cpu.rf_ram.memory[264][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[265][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[266][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[267][1] ),
    .S0(_01802_),
    .S1(_01932_),
    .Z(_02899_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08593_ (.A1(_01979_),
    .A2(_02899_),
    .B(_01788_),
    .ZN(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08594_ (.I0(\mod.u_cpu.rf_ram.memory[256][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[257][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[258][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[259][1] ),
    .S0(_01837_),
    .S1(_02252_),
    .Z(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08595_ (.I(\mod.u_cpu.rf_ram.memory[261][1] ),
    .ZN(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08596_ (.A1(_01858_),
    .A2(_02902_),
    .ZN(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08597_ (.A1(_02070_),
    .A2(\mod.u_cpu.rf_ram.memory[260][1] ),
    .B(_02903_),
    .ZN(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08598_ (.I(\mod.u_cpu.rf_ram.memory[263][1] ),
    .ZN(_02905_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08599_ (.A1(_01672_),
    .A2(_02905_),
    .ZN(_02906_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08600_ (.A1(_02136_),
    .A2(\mod.u_cpu.rf_ram.memory[262][1] ),
    .B(_02906_),
    .C(_01504_),
    .ZN(_02907_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08601_ (.A1(_02323_),
    .A2(_02904_),
    .B(_02907_),
    .C(_01631_),
    .ZN(_02908_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08602_ (.A1(_01852_),
    .A2(_02901_),
    .B(_02908_),
    .C(_01887_),
    .ZN(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08603_ (.A1(_02898_),
    .A2(_02900_),
    .B(_02046_),
    .C(_02909_),
    .ZN(_02910_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08604_ (.A1(_01977_),
    .A2(_02893_),
    .A3(_02910_),
    .ZN(_02911_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08605_ (.A1(_01738_),
    .A2(_02874_),
    .A3(_02911_),
    .ZN(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08606_ (.A1(_01470_),
    .A2(_02836_),
    .A3(_02912_),
    .Z(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08607_ (.A1(_01481_),
    .A2(_02758_),
    .B(_02913_),
    .C(_01469_),
    .ZN(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08608_ (.I0(\mod.u_cpu.rf_ram.memory[128][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[129][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[130][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[131][1] ),
    .S0(_02638_),
    .S1(_02067_),
    .Z(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08609_ (.A1(_02040_),
    .A2(_02915_),
    .ZN(_02916_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08610_ (.I0(\mod.u_cpu.rf_ram.memory[144][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[145][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[146][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[147][1] ),
    .S0(_02085_),
    .S1(_02049_),
    .Z(_02917_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08611_ (.A1(_02074_),
    .A2(_02917_),
    .B(_01662_),
    .ZN(_02918_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08612_ (.I0(\mod.u_cpu.rf_ram.memory[132][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[133][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[134][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[135][1] ),
    .S0(_01893_),
    .S1(_02054_),
    .Z(_02919_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08613_ (.A1(_02053_),
    .A2(_02919_),
    .ZN(_02920_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08614_ (.I0(\mod.u_cpu.rf_ram.memory[148][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[149][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[150][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[151][1] ),
    .S0(_02059_),
    .S1(_01723_),
    .Z(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08615_ (.A1(_02057_),
    .A2(_02921_),
    .B(_01632_),
    .ZN(_02922_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08616_ (.A1(_02916_),
    .A2(_02918_),
    .B1(_02920_),
    .B2(_02922_),
    .C(_01658_),
    .ZN(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08617_ (.I0(\mod.u_cpu.rf_ram.memory[136][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[137][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[138][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[139][1] ),
    .S0(_02022_),
    .S1(_02043_),
    .Z(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08618_ (.A1(_01849_),
    .A2(_02924_),
    .ZN(_02925_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08619_ (.I0(\mod.u_cpu.rf_ram.memory[152][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[153][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[154][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[155][1] ),
    .S0(_02066_),
    .S1(_02067_),
    .Z(_02926_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08620_ (.A1(_02046_),
    .A2(_02926_),
    .B(_02051_),
    .ZN(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08621_ (.I0(\mod.u_cpu.rf_ram.memory[140][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[141][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[142][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[143][1] ),
    .S0(_02070_),
    .S1(_02071_),
    .Z(_02928_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08622_ (.A1(_02053_),
    .A2(_02928_),
    .ZN(_02929_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08623_ (.I0(\mod.u_cpu.rf_ram.memory[156][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[157][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[158][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[159][1] ),
    .S0(_01925_),
    .S1(_02071_),
    .Z(_02930_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08624_ (.A1(_02074_),
    .A2(_02930_),
    .B(_01602_),
    .ZN(_02931_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08625_ (.A1(_02925_),
    .A2(_02927_),
    .B1(_02929_),
    .B2(_02931_),
    .C(_02077_),
    .ZN(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08626_ (.A1(_01486_),
    .A2(_02923_),
    .A3(_02932_),
    .Z(_02933_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08627_ (.I0(\mod.u_cpu.rf_ram.memory[176][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[177][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[178][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[179][1] ),
    .S0(_02048_),
    .S1(_02086_),
    .Z(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08628_ (.A1(_02090_),
    .A2(_02934_),
    .ZN(_02935_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08629_ (.I0(\mod.u_cpu.rf_ram.memory[180][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[181][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[182][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[183][1] ),
    .S0(_02085_),
    .S1(_02086_),
    .Z(_02936_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08630_ (.A1(_02097_),
    .A2(_02936_),
    .ZN(_02937_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08631_ (.A1(_01818_),
    .A2(_02935_),
    .A3(_02937_),
    .ZN(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08632_ (.I0(\mod.u_cpu.rf_ram.memory[184][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[185][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[186][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[187][1] ),
    .S0(_02092_),
    .S1(_02098_),
    .Z(_02939_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08633_ (.A1(_02090_),
    .A2(_02939_),
    .ZN(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08634_ (.I0(\mod.u_cpu.rf_ram.memory[188][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[189][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[190][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[191][1] ),
    .S0(_02092_),
    .S1(_02098_),
    .Z(_02941_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08635_ (.A1(_02097_),
    .A2(_02941_),
    .ZN(_02942_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08636_ (.A1(_01836_),
    .A2(_02940_),
    .A3(_02942_),
    .ZN(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08637_ (.A1(_02938_),
    .A2(_02943_),
    .B(_02102_),
    .ZN(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08638_ (.I0(\mod.u_cpu.rf_ram.memory[168][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[169][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[170][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[171][1] ),
    .S0(_02106_),
    .S1(_02127_),
    .Z(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08639_ (.I(\mod.u_cpu.rf_ram.memory[173][1] ),
    .ZN(_02946_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08640_ (.A1(_02130_),
    .A2(_02946_),
    .ZN(_02947_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08641_ (.A1(_02111_),
    .A2(\mod.u_cpu.rf_ram.memory[172][1] ),
    .B(_02947_),
    .ZN(_02948_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08642_ (.I(\mod.u_cpu.rf_ram.memory[175][1] ),
    .ZN(_02949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08643_ (.A1(_02116_),
    .A2(_02949_),
    .ZN(_02950_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08644_ (.A1(_02115_),
    .A2(\mod.u_cpu.rf_ram.memory[174][1] ),
    .B(_02950_),
    .C(_01771_),
    .ZN(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08645_ (.A1(_02110_),
    .A2(_02948_),
    .B(_02951_),
    .C(_02141_),
    .ZN(_02952_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08646_ (.A1(_01670_),
    .A2(_02945_),
    .B(_02952_),
    .C(_02122_),
    .ZN(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08647_ (.I0(\mod.u_cpu.rf_ram.memory[160][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[161][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[162][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[163][1] ),
    .S0(_02125_),
    .S1(_02127_),
    .Z(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08648_ (.I(\mod.u_cpu.rf_ram.memory[165][1] ),
    .ZN(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08649_ (.A1(_02130_),
    .A2(_02955_),
    .ZN(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08650_ (.A1(_02129_),
    .A2(\mod.u_cpu.rf_ram.memory[164][1] ),
    .B(_02956_),
    .ZN(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08651_ (.I(\mod.u_cpu.rf_ram.memory[167][1] ),
    .ZN(_02958_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08652_ (.A1(_02136_),
    .A2(_02958_),
    .ZN(_02959_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08653_ (.A1(_02135_),
    .A2(\mod.u_cpu.rf_ram.memory[166][1] ),
    .B(_02959_),
    .C(_02139_),
    .ZN(_02960_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08654_ (.A1(_02110_),
    .A2(_02957_),
    .B(_02960_),
    .C(_02141_),
    .ZN(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08655_ (.A1(_02124_),
    .A2(_02954_),
    .B(_02961_),
    .C(_02143_),
    .ZN(_02962_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08656_ (.A1(_02105_),
    .A2(_02953_),
    .A3(_02962_),
    .ZN(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08657_ (.A1(_02104_),
    .A2(_02963_),
    .ZN(_02964_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08658_ (.A1(_02944_),
    .A2(_02964_),
    .B(_01738_),
    .ZN(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08659_ (.I(\mod.u_cpu.rf_ram.memory[221][1] ),
    .ZN(_02966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08660_ (.A1(_02656_),
    .A2(_02966_),
    .ZN(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08661_ (.A1(_02450_),
    .A2(\mod.u_cpu.rf_ram.memory[220][1] ),
    .B(_02967_),
    .ZN(_02968_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08662_ (.I(\mod.u_cpu.rf_ram.memory[223][1] ),
    .ZN(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08663_ (.A1(_02711_),
    .A2(_02969_),
    .ZN(_02970_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08664_ (.A1(_02566_),
    .A2(\mod.u_cpu.rf_ram.memory[222][1] ),
    .B(_02970_),
    .C(_01703_),
    .ZN(_02971_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08665_ (.A1(_02561_),
    .A2(_02968_),
    .B(_02971_),
    .C(_01696_),
    .ZN(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08666_ (.I0(\mod.u_cpu.rf_ram.memory[218][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[219][1] ),
    .S(_02294_),
    .Z(_02973_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08667_ (.I(\mod.u_cpu.rf_ram.memory[217][1] ),
    .ZN(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08668_ (.A1(_01567_),
    .A2(\mod.u_cpu.rf_ram.memory[216][1] ),
    .ZN(_02975_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08669_ (.A1(_02711_),
    .A2(_02974_),
    .B(_02975_),
    .C(_01723_),
    .ZN(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08670_ (.A1(_02759_),
    .A2(_02973_),
    .B(_02976_),
    .C(_01872_),
    .ZN(_02977_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08671_ (.A1(_02606_),
    .A2(_02977_),
    .ZN(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08672_ (.I(\mod.u_cpu.rf_ram.memory[213][1] ),
    .ZN(_02979_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08673_ (.A1(_02202_),
    .A2(_02979_),
    .ZN(_02980_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08674_ (.A1(_02479_),
    .A2(\mod.u_cpu.rf_ram.memory[212][1] ),
    .B(_02980_),
    .ZN(_02981_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08675_ (.I(\mod.u_cpu.rf_ram.memory[215][1] ),
    .ZN(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08676_ (.A1(_01705_),
    .A2(_02982_),
    .ZN(_02983_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08677_ (.A1(_02462_),
    .A2(\mod.u_cpu.rf_ram.memory[214][1] ),
    .B(_02983_),
    .C(_02597_),
    .ZN(_02984_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08678_ (.A1(_02543_),
    .A2(_02981_),
    .B(_02984_),
    .C(_01632_),
    .ZN(_02985_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08679_ (.I0(\mod.u_cpu.rf_ram.memory[210][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[211][1] ),
    .S(_01807_),
    .Z(_02986_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08680_ (.I(\mod.u_cpu.rf_ram.memory[209][1] ),
    .ZN(_02987_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08681_ (.A1(_02632_),
    .A2(\mod.u_cpu.rf_ram.memory[208][1] ),
    .ZN(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08682_ (.A1(_02477_),
    .A2(_02987_),
    .B(_02988_),
    .C(_01638_),
    .ZN(_02989_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08683_ (.A1(_02594_),
    .A2(_02986_),
    .B(_02989_),
    .C(_02591_),
    .ZN(_02990_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08684_ (.A1(_02230_),
    .A2(_02990_),
    .ZN(_02991_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08685_ (.A1(_02972_),
    .A2(_02978_),
    .B1(_02985_),
    .B2(_02991_),
    .C(_01489_),
    .ZN(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08686_ (.I0(\mod.u_cpu.rf_ram.memory[206][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[207][1] ),
    .S(_01545_),
    .Z(_02993_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08687_ (.I(\mod.u_cpu.rf_ram.memory[205][1] ),
    .ZN(_02994_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08688_ (.A1(_02179_),
    .A2(\mod.u_cpu.rf_ram.memory[204][1] ),
    .ZN(_02995_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08689_ (.A1(_02202_),
    .A2(_02994_),
    .B(_02995_),
    .C(_02093_),
    .ZN(_02996_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08690_ (.A1(_02578_),
    .A2(_02993_),
    .B(_02996_),
    .C(_02660_),
    .ZN(_02997_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08691_ (.I0(\mod.u_cpu.rf_ram.memory[200][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[201][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[202][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[203][1] ),
    .S0(_02349_),
    .S1(_02350_),
    .Z(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08692_ (.A1(_02348_),
    .A2(_02998_),
    .B(_02377_),
    .ZN(_02999_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08693_ (.I0(\mod.u_cpu.rf_ram.memory[192][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[193][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[194][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[195][1] ),
    .S0(_01578_),
    .S1(_01714_),
    .Z(_03000_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08694_ (.I(_01560_),
    .Z(_03001_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08695_ (.I(\mod.u_cpu.rf_ram.memory[197][1] ),
    .ZN(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08696_ (.A1(_03001_),
    .A2(_03002_),
    .ZN(_03003_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08697_ (.A1(_02204_),
    .A2(\mod.u_cpu.rf_ram.memory[196][1] ),
    .B(_03003_),
    .ZN(_03004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08698_ (.I(\mod.u_cpu.rf_ram.memory[199][1] ),
    .ZN(_03005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08699_ (.A1(_02190_),
    .A2(_03005_),
    .ZN(_03006_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08700_ (.A1(_01573_),
    .A2(\mod.u_cpu.rf_ram.memory[198][1] ),
    .B(_03006_),
    .C(_02212_),
    .ZN(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08701_ (.A1(_02063_),
    .A2(_03004_),
    .B(_03007_),
    .C(_01669_),
    .ZN(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08702_ (.A1(_02665_),
    .A2(_03000_),
    .B(_03008_),
    .C(_02852_),
    .ZN(_03009_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08703_ (.A1(_02997_),
    .A2(_02999_),
    .B(_01891_),
    .C(_03009_),
    .ZN(_03010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08704_ (.A1(_01486_),
    .A2(_03010_),
    .ZN(_03011_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08705_ (.I0(\mod.u_cpu.rf_ram.memory[238][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[239][1] ),
    .S(_01807_),
    .Z(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08706_ (.I(\mod.u_cpu.rf_ram.memory[237][1] ),
    .ZN(_03013_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08707_ (.A1(_02385_),
    .A2(\mod.u_cpu.rf_ram.memory[236][1] ),
    .ZN(_03014_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08708_ (.A1(_02209_),
    .A2(_03013_),
    .B(_03014_),
    .C(_02633_),
    .ZN(_03015_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08709_ (.A1(_02594_),
    .A2(_03012_),
    .B(_03015_),
    .C(_02764_),
    .ZN(_03016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08710_ (.I(_01991_),
    .Z(_03017_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08711_ (.I0(\mod.u_cpu.rf_ram.memory[232][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[233][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[234][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[235][1] ),
    .S0(_01647_),
    .S1(_01732_),
    .Z(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08712_ (.A1(_03017_),
    .A2(_03018_),
    .B(_01870_),
    .ZN(_03019_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08713_ (.I0(\mod.u_cpu.rf_ram.memory[224][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[225][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[226][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[227][1] ),
    .S0(_01507_),
    .S1(_01763_),
    .Z(_03020_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08714_ (.I(\mod.u_cpu.rf_ram.memory[229][1] ),
    .ZN(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08715_ (.A1(_02027_),
    .A2(_03021_),
    .ZN(_03022_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08716_ (.A1(_01608_),
    .A2(\mod.u_cpu.rf_ram.memory[228][1] ),
    .B(_03022_),
    .ZN(_03023_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08717_ (.I(\mod.u_cpu.rf_ram.memory[231][1] ),
    .ZN(_03024_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08718_ (.A1(_01704_),
    .A2(_03024_),
    .ZN(_03025_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08719_ (.A1(_02751_),
    .A2(\mod.u_cpu.rf_ram.memory[230][1] ),
    .B(_03025_),
    .C(_02154_),
    .ZN(_03026_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08720_ (.A1(_01698_),
    .A2(_03023_),
    .B(_03026_),
    .C(_02347_),
    .ZN(_03027_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08721_ (.A1(_02591_),
    .A2(_03020_),
    .B(_03027_),
    .C(_01657_),
    .ZN(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08722_ (.A1(_03016_),
    .A2(_03019_),
    .B(_02074_),
    .C(_03028_),
    .ZN(_03029_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08723_ (.I0(\mod.u_cpu.rf_ram.memory[240][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[241][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[242][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[243][1] ),
    .S0(_01647_),
    .S1(_01732_),
    .Z(_03030_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08724_ (.I(\mod.u_cpu.rf_ram.memory[245][1] ),
    .ZN(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08725_ (.A1(_02197_),
    .A2(_03031_),
    .ZN(_03032_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08726_ (.A1(_02161_),
    .A2(\mod.u_cpu.rf_ram.memory[244][1] ),
    .B(_03032_),
    .ZN(_03033_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08727_ (.I(\mod.u_cpu.rf_ram.memory[247][1] ),
    .ZN(_03034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08728_ (.A1(_02084_),
    .A2(_03034_),
    .ZN(_03035_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08729_ (.A1(_02632_),
    .A2(\mod.u_cpu.rf_ram.memory[246][1] ),
    .B(_03035_),
    .C(_01702_),
    .ZN(_03036_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08730_ (.A1(_02043_),
    .A2(_03033_),
    .B(_03036_),
    .C(_01695_),
    .ZN(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08731_ (.A1(_03017_),
    .A2(_03030_),
    .B(_03037_),
    .C(_02852_),
    .ZN(_03038_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08732_ (.I0(\mod.u_cpu.rf_ram.memory[248][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[249][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[250][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[251][1] ),
    .S0(_03001_),
    .S1(_01525_),
    .Z(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08733_ (.I(\mod.u_cpu.rf_ram.memory[253][1] ),
    .ZN(_03040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08734_ (.A1(_02197_),
    .A2(_03040_),
    .ZN(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08735_ (.A1(_02179_),
    .A2(\mod.u_cpu.rf_ram.memory[252][1] ),
    .B(_03041_),
    .ZN(_03042_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08736_ (.I(\mod.u_cpu.rf_ram.memory[255][1] ),
    .ZN(_03043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08737_ (.A1(_02084_),
    .A2(_03043_),
    .ZN(_03044_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08738_ (.A1(_02632_),
    .A2(\mod.u_cpu.rf_ram.memory[254][1] ),
    .B(_03044_),
    .C(_01702_),
    .ZN(_03045_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08739_ (.A1(_02043_),
    .A2(_03042_),
    .B(_03045_),
    .C(_01695_),
    .ZN(_03046_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08740_ (.A1(_03017_),
    .A2(_03039_),
    .B(_03046_),
    .C(_01870_),
    .ZN(_03047_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08741_ (.A1(_01978_),
    .A2(_03038_),
    .A3(_03047_),
    .ZN(_03048_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08742_ (.A1(_01848_),
    .A2(_03029_),
    .A3(_03048_),
    .ZN(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08743_ (.A1(_02992_),
    .A2(_03011_),
    .B(_03049_),
    .C(_02148_),
    .ZN(_03050_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08744_ (.A1(_02933_),
    .A2(_02965_),
    .B(_01481_),
    .C(_03050_),
    .ZN(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08745_ (.I0(\mod.u_cpu.rf_ram.memory[110][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[111][1] ),
    .S(_01508_),
    .Z(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08746_ (.I(\mod.u_cpu.rf_ram.memory[109][1] ),
    .ZN(_03053_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08747_ (.A1(_02156_),
    .A2(\mod.u_cpu.rf_ram.memory[108][1] ),
    .ZN(_03054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08748_ (.A1(_02585_),
    .A2(_03053_),
    .B(_03054_),
    .C(_01751_),
    .ZN(_03055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08749_ (.A1(_02611_),
    .A2(_03052_),
    .B(_03055_),
    .C(_01680_),
    .ZN(_03056_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08750_ (.I0(\mod.u_cpu.rf_ram.memory[104][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[105][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[106][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[107][1] ),
    .S0(_02106_),
    .S1(_02107_),
    .Z(_03057_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08751_ (.A1(_01670_),
    .A2(_03057_),
    .B(_02230_),
    .ZN(_03058_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08752_ (.I0(\mod.u_cpu.rf_ram.memory[96][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[97][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[98][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[99][1] ),
    .S0(_02211_),
    .S1(_02386_),
    .Z(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08753_ (.I(\mod.u_cpu.rf_ram.memory[101][1] ),
    .ZN(_03060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08754_ (.A1(_02171_),
    .A2(_03060_),
    .ZN(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08755_ (.A1(_02532_),
    .A2(\mod.u_cpu.rf_ram.memory[100][1] ),
    .B(_03061_),
    .ZN(_03062_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08756_ (.I(\mod.u_cpu.rf_ram.memory[103][1] ),
    .ZN(_03063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08757_ (.A1(_02220_),
    .A2(_03063_),
    .ZN(_03064_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08758_ (.A1(_02204_),
    .A2(\mod.u_cpu.rf_ram.memory[102][1] ),
    .B(_03064_),
    .C(_02359_),
    .ZN(_03065_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08759_ (.A1(_02352_),
    .A2(_03062_),
    .B(_03065_),
    .C(_02361_),
    .ZN(_03066_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08760_ (.A1(_02631_),
    .A2(_03059_),
    .B(_03066_),
    .C(_02363_),
    .ZN(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08761_ (.A1(_03056_),
    .A2(_03058_),
    .B(_02149_),
    .C(_03067_),
    .ZN(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08762_ (.I0(\mod.u_cpu.rf_ram.memory[120][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[121][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[122][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[123][1] ),
    .S0(_02294_),
    .S1(_02295_),
    .Z(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08763_ (.I(\mod.u_cpu.rf_ram.memory[125][1] ),
    .ZN(_03070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08764_ (.A1(_02298_),
    .A2(_03070_),
    .ZN(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08765_ (.A1(_02297_),
    .A2(\mod.u_cpu.rf_ram.memory[124][1] ),
    .B(_03071_),
    .ZN(_03072_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08766_ (.I(\mod.u_cpu.rf_ram.memory[127][1] ),
    .ZN(_03073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08767_ (.A1(_02303_),
    .A2(_03073_),
    .ZN(_03074_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08768_ (.A1(_02316_),
    .A2(\mod.u_cpu.rf_ram.memory[126][1] ),
    .B(_03074_),
    .C(_02306_),
    .ZN(_03075_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08769_ (.A1(_02283_),
    .A2(_03072_),
    .B(_03075_),
    .C(_02308_),
    .ZN(_03076_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08770_ (.A1(_02293_),
    .A2(_03069_),
    .B(_03076_),
    .C(_02321_),
    .ZN(_03077_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08771_ (.I0(\mod.u_cpu.rf_ram.memory[112][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[113][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[114][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[115][1] ),
    .S0(_01664_),
    .S1(_02323_),
    .Z(_03078_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08772_ (.I(\mod.u_cpu.rf_ram.memory[117][1] ),
    .ZN(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08773_ (.A1(_01682_),
    .A2(_03079_),
    .ZN(_03080_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08774_ (.A1(_02477_),
    .A2(\mod.u_cpu.rf_ram.memory[116][1] ),
    .B(_03080_),
    .ZN(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08775_ (.I(\mod.u_cpu.rf_ram.memory[119][1] ),
    .ZN(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08776_ (.A1(_01863_),
    .A2(_03082_),
    .ZN(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08777_ (.A1(_02329_),
    .A2(\mod.u_cpu.rf_ram.memory[118][1] ),
    .B(_03083_),
    .C(_01916_),
    .ZN(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08778_ (.A1(_02325_),
    .A2(_03081_),
    .B(_03084_),
    .C(_01717_),
    .ZN(_03085_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08779_ (.A1(_01688_),
    .A2(_03078_),
    .B(_03085_),
    .C(_02291_),
    .ZN(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08780_ (.A1(_01446_),
    .A2(_03077_),
    .A3(_03086_),
    .ZN(_03087_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08781_ (.A1(_02104_),
    .A2(_03068_),
    .A3(_03087_),
    .ZN(_03088_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08782_ (.I0(\mod.u_cpu.rf_ram.memory[80][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[81][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[82][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[83][1] ),
    .S0(_02249_),
    .S1(_02107_),
    .Z(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08783_ (.A1(_02051_),
    .A2(_03089_),
    .ZN(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08784_ (.I0(\mod.u_cpu.rf_ram.memory[84][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[85][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[86][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[87][1] ),
    .S0(_01857_),
    .S1(_02054_),
    .Z(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08785_ (.A1(_01696_),
    .A2(_03091_),
    .B(_01720_),
    .ZN(_03092_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08786_ (.I0(\mod.u_cpu.rf_ram.memory[88][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[89][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[90][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[91][1] ),
    .S0(_01673_),
    .S1(_01855_),
    .Z(_03093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08787_ (.A1(_01662_),
    .A2(_03093_),
    .ZN(_03094_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08788_ (.I0(\mod.u_cpu.rf_ram.memory[92][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[93][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[94][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[95][1] ),
    .S0(_01636_),
    .S1(_01638_),
    .Z(_03095_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08789_ (.A1(_01493_),
    .A2(_03095_),
    .B(_01534_),
    .ZN(_03096_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08790_ (.A1(_03090_),
    .A2(_03092_),
    .B1(_03094_),
    .B2(_03096_),
    .ZN(_03097_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08791_ (.I0(\mod.u_cpu.rf_ram.memory[78][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[79][1] ),
    .S(_01517_),
    .Z(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08792_ (.I(\mod.u_cpu.rf_ram.memory[77][1] ),
    .ZN(_03099_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08793_ (.A1(_02161_),
    .A2(\mod.u_cpu.rf_ram.memory[76][1] ),
    .ZN(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08794_ (.A1(_02202_),
    .A2(_03099_),
    .B(_03100_),
    .C(_02086_),
    .ZN(_03101_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08795_ (.A1(_02465_),
    .A2(_03098_),
    .B(_03101_),
    .C(_02660_),
    .ZN(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08796_ (.I0(\mod.u_cpu.rf_ram.memory[72][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[73][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[74][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[75][1] ),
    .S0(_02211_),
    .S1(_02386_),
    .Z(_03103_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08797_ (.A1(_02348_),
    .A2(_03103_),
    .B(_01618_),
    .ZN(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08798_ (.I0(\mod.u_cpu.rf_ram.memory[64][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[65][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[66][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[67][1] ),
    .S0(_01561_),
    .S1(_01714_),
    .Z(_03105_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08799_ (.I(\mod.u_cpu.rf_ram.memory[69][1] ),
    .ZN(_03106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08800_ (.A1(_03001_),
    .A2(_03106_),
    .ZN(_03107_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08801_ (.A1(_02204_),
    .A2(\mod.u_cpu.rf_ram.memory[68][1] ),
    .B(_03107_),
    .ZN(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08802_ (.I(\mod.u_cpu.rf_ram.memory[71][1] ),
    .ZN(_03109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08803_ (.A1(_02190_),
    .A2(_03109_),
    .ZN(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08804_ (.A1(_01511_),
    .A2(\mod.u_cpu.rf_ram.memory[70][1] ),
    .B(_03110_),
    .C(_02109_),
    .ZN(_03111_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08805_ (.A1(_02063_),
    .A2(_03108_),
    .B(_03111_),
    .C(_01669_),
    .ZN(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08806_ (.A1(_02665_),
    .A2(_03105_),
    .B(_03112_),
    .C(_02677_),
    .ZN(_03113_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08807_ (.A1(_03102_),
    .A2(_03104_),
    .B(_03113_),
    .C(_02664_),
    .ZN(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08808_ (.A1(_02337_),
    .A2(_03097_),
    .B(_03114_),
    .C(_02380_),
    .ZN(_03115_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08809_ (.A1(_01483_),
    .A2(_03088_),
    .A3(_03115_),
    .ZN(_03116_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08810_ (.I0(\mod.u_cpu.rf_ram.memory[4][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[5][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[6][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[7][1] ),
    .S0(_02366_),
    .S1(_02383_),
    .Z(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08811_ (.I0(\mod.u_cpu.rf_ram.memory[0][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[1][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[2][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[3][1] ),
    .S0(_02211_),
    .S1(_02386_),
    .Z(_03118_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08812_ (.I0(\mod.u_cpu.rf_ram.memory[12][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[13][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[14][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[15][1] ),
    .S0(_02266_),
    .S1(_02388_),
    .Z(_03119_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08813_ (.I0(\mod.u_cpu.rf_ram.memory[8][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[9][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[10][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[11][1] ),
    .S0(_02171_),
    .S1(_02267_),
    .Z(_03120_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08814_ (.I0(_03117_),
    .I1(_03118_),
    .I2(_03119_),
    .I3(_03120_),
    .S0(_02391_),
    .S1(_01720_),
    .Z(_03121_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08815_ (.I0(\mod.u_cpu.rf_ram.memory[24][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[25][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[26][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[27][1] ),
    .S0(_02366_),
    .S1(_02367_),
    .Z(_03122_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08816_ (.I(\mod.u_cpu.rf_ram.memory[29][1] ),
    .ZN(_03123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08817_ (.A1(_02369_),
    .A2(_03123_),
    .ZN(_03124_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08818_ (.A1(_02302_),
    .A2(\mod.u_cpu.rf_ram.memory[28][1] ),
    .B(_03124_),
    .ZN(_03125_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08819_ (.I(\mod.u_cpu.rf_ram.memory[31][1] ),
    .ZN(_03126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08820_ (.A1(_02411_),
    .A2(_03126_),
    .ZN(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08821_ (.A1(_02410_),
    .A2(\mod.u_cpu.rf_ram.memory[30][1] ),
    .B(_03127_),
    .C(_01830_),
    .ZN(_03128_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08822_ (.A1(_02405_),
    .A2(_03125_),
    .B(_03128_),
    .C(_02415_),
    .ZN(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08823_ (.A1(_02365_),
    .A2(_03122_),
    .B(_03129_),
    .C(_02185_),
    .ZN(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08824_ (.I0(\mod.u_cpu.rf_ram.memory[16][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[17][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[18][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[19][1] ),
    .S0(_02403_),
    .S1(_02367_),
    .Z(_03131_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08825_ (.I(\mod.u_cpu.rf_ram.memory[21][1] ),
    .ZN(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08826_ (.A1(_02406_),
    .A2(_03132_),
    .ZN(_03133_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08827_ (.A1(_02316_),
    .A2(\mod.u_cpu.rf_ram.memory[20][1] ),
    .B(_03133_),
    .ZN(_03134_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08828_ (.I(\mod.u_cpu.rf_ram.memory[23][1] ),
    .ZN(_03135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08829_ (.A1(_02411_),
    .A2(_03135_),
    .ZN(_03136_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08830_ (.A1(_02410_),
    .A2(\mod.u_cpu.rf_ram.memory[22][1] ),
    .B(_03136_),
    .C(_01830_),
    .ZN(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08831_ (.A1(_02405_),
    .A2(_03134_),
    .B(_03137_),
    .C(_02415_),
    .ZN(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08832_ (.A1(_02150_),
    .A2(_03131_),
    .B(_03138_),
    .C(_02363_),
    .ZN(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08833_ (.A1(_01592_),
    .A2(_03130_),
    .A3(_03139_),
    .ZN(_03140_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08834_ (.A1(_01693_),
    .A2(_03121_),
    .B(_03140_),
    .C(_02380_),
    .ZN(_03141_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08835_ (.I0(\mod.u_cpu.rf_ram.memory[52][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[53][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[54][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[55][1] ),
    .S0(_02151_),
    .S1(_02152_),
    .Z(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08836_ (.I0(\mod.u_cpu.rf_ram.memory[48][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[49][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[50][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[51][1] ),
    .S0(_02421_),
    .S1(_02393_),
    .Z(_03143_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08837_ (.I0(\mod.u_cpu.rf_ram.memory[60][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[61][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[62][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[63][1] ),
    .S0(_02406_),
    .S1(_02218_),
    .Z(_03144_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08838_ (.I0(\mod.u_cpu.rf_ram.memory[56][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[57][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[58][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[59][1] ),
    .S0(_02242_),
    .S1(_02388_),
    .Z(_03145_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08839_ (.I0(_03142_),
    .I1(_03143_),
    .I2(_03144_),
    .I3(_03145_),
    .S0(_02391_),
    .S1(_01552_),
    .Z(_03146_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08840_ (.I0(\mod.u_cpu.rf_ram.memory[46][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[47][1] ),
    .S(_01577_),
    .Z(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08841_ (.I(\mod.u_cpu.rf_ram.memory[45][1] ),
    .ZN(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08842_ (.A1(_02272_),
    .A2(\mod.u_cpu.rf_ram.memory[44][1] ),
    .ZN(_03149_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08843_ (.A1(_02191_),
    .A2(_03148_),
    .B(_03149_),
    .C(_02093_),
    .ZN(_03150_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08844_ (.A1(_02578_),
    .A2(_03147_),
    .B(_03150_),
    .C(_02660_),
    .ZN(_03151_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08845_ (.I0(\mod.u_cpu.rf_ram.memory[40][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[41][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[42][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[43][1] ),
    .S0(_02349_),
    .S1(_02393_),
    .Z(_03152_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08846_ (.A1(_02365_),
    .A2(_03152_),
    .B(_02377_),
    .ZN(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08847_ (.I0(\mod.u_cpu.rf_ram.memory[32][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[33][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[34][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[35][1] ),
    .S0(_01647_),
    .S1(_01732_),
    .Z(_03154_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08848_ (.I(\mod.u_cpu.rf_ram.memory[37][1] ),
    .ZN(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08849_ (.A1(_03001_),
    .A2(_03155_),
    .ZN(_03156_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08850_ (.A1(_02356_),
    .A2(\mod.u_cpu.rf_ram.memory[36][1] ),
    .B(_03156_),
    .ZN(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08851_ (.I(\mod.u_cpu.rf_ram.memory[39][1] ),
    .ZN(_03158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08852_ (.A1(_02190_),
    .A2(_03158_),
    .ZN(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08853_ (.A1(_01608_),
    .A2(\mod.u_cpu.rf_ram.memory[38][1] ),
    .B(_03159_),
    .C(_02212_),
    .ZN(_03160_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08854_ (.A1(_02063_),
    .A2(_03157_),
    .B(_03160_),
    .C(_01695_),
    .ZN(_03161_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08855_ (.A1(_03017_),
    .A2(_03154_),
    .B(_03161_),
    .C(_02852_),
    .ZN(_03162_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08856_ (.A1(_03151_),
    .A2(_03153_),
    .B(_03162_),
    .C(_01891_),
    .ZN(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08857_ (.A1(_02102_),
    .A2(_03146_),
    .B(_03163_),
    .C(_01739_),
    .ZN(_03164_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08858_ (.A1(_01475_),
    .A2(_03141_),
    .A3(_03164_),
    .ZN(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08859_ (.A1(_01471_),
    .A2(_03116_),
    .A3(_03165_),
    .ZN(_03166_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08860_ (.A1(_01468_),
    .A2(_03051_),
    .A3(_03166_),
    .Z(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08861_ (.I0(\mod.u_cpu.rf_ram.memory[544][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[545][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[546][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[547][1] ),
    .S0(_02450_),
    .S1(_02451_),
    .Z(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08862_ (.I(\mod.u_cpu.rf_ram.memory[549][1] ),
    .ZN(_03169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08863_ (.A1(_02472_),
    .A2(_03169_),
    .ZN(_03170_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08864_ (.A1(_02456_),
    .A2(\mod.u_cpu.rf_ram.memory[548][1] ),
    .B(_03170_),
    .ZN(_03171_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08865_ (.I(\mod.u_cpu.rf_ram.memory[551][1] ),
    .ZN(_03172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08866_ (.A1(_02462_),
    .A2(_03172_),
    .ZN(_03173_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08867_ (.A1(_02461_),
    .A2(\mod.u_cpu.rf_ram.memory[550][1] ),
    .B(_03173_),
    .C(_02578_),
    .ZN(_03174_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08868_ (.A1(_02455_),
    .A2(_03171_),
    .B(_03174_),
    .C(_02555_),
    .ZN(_03175_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08869_ (.A1(_02542_),
    .A2(_03168_),
    .B(_03175_),
    .C(_02518_),
    .ZN(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08870_ (.I0(\mod.u_cpu.rf_ram.memory[552][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[553][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[554][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[555][1] ),
    .S0(_02472_),
    .S1(_02473_),
    .Z(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08871_ (.I(\mod.u_cpu.rf_ram.memory[557][1] ),
    .ZN(_03178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08872_ (.A1(_02479_),
    .A2(_03178_),
    .ZN(_03179_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08873_ (.A1(_02478_),
    .A2(\mod.u_cpu.rf_ram.memory[556][1] ),
    .B(_03179_),
    .ZN(_03180_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08874_ (.I(\mod.u_cpu.rf_ram.memory[559][1] ),
    .ZN(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08875_ (.A1(_02484_),
    .A2(_03181_),
    .ZN(_03182_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08876_ (.A1(_02483_),
    .A2(\mod.u_cpu.rf_ram.memory[558][1] ),
    .B(_03182_),
    .C(_02487_),
    .ZN(_03183_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08877_ (.A1(_02476_),
    .A2(_03180_),
    .B(_03183_),
    .C(_02083_),
    .ZN(_03184_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08878_ (.A1(_02592_),
    .A2(_03177_),
    .B(_03184_),
    .C(_01836_),
    .ZN(_03185_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08879_ (.A1(_03176_),
    .A2(_03185_),
    .B(_02609_),
    .ZN(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08880_ (.I0(\mod.u_cpu.rf_ram.memory[568][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[569][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[570][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[571][1] ),
    .S0(_02494_),
    .S1(_02451_),
    .Z(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08881_ (.I(\mod.u_cpu.rf_ram.memory[573][1] ),
    .ZN(_03188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08882_ (.A1(_02457_),
    .A2(_03188_),
    .ZN(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08883_ (.A1(_02456_),
    .A2(\mod.u_cpu.rf_ram.memory[572][1] ),
    .B(_03189_),
    .ZN(_03190_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08884_ (.I(\mod.u_cpu.rf_ram.memory[575][1] ),
    .ZN(_03191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08885_ (.A1(_02500_),
    .A2(_03191_),
    .ZN(_03192_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08886_ (.A1(_02461_),
    .A2(\mod.u_cpu.rf_ram.memory[574][1] ),
    .B(_03192_),
    .C(_02465_),
    .ZN(_03193_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08887_ (.A1(_02455_),
    .A2(_03190_),
    .B(_03193_),
    .C(_02467_),
    .ZN(_03194_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08888_ (.A1(_02449_),
    .A2(_03187_),
    .B(_03194_),
    .C(_02505_),
    .ZN(_03195_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08889_ (.I0(\mod.u_cpu.rf_ram.memory[560][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[561][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[562][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[563][1] ),
    .S0(_02457_),
    .S1(_02473_),
    .Z(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08890_ (.I(\mod.u_cpu.rf_ram.memory[565][1] ),
    .ZN(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08891_ (.A1(_02479_),
    .A2(_03197_),
    .ZN(_03198_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08892_ (.A1(_02478_),
    .A2(\mod.u_cpu.rf_ram.memory[564][1] ),
    .B(_03198_),
    .ZN(_03199_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08893_ (.I(\mod.u_cpu.rf_ram.memory[567][1] ),
    .ZN(_03200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08894_ (.A1(_02484_),
    .A2(_03200_),
    .ZN(_03201_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08895_ (.A1(_02483_),
    .A2(\mod.u_cpu.rf_ram.memory[566][1] ),
    .B(_03201_),
    .C(_02487_),
    .ZN(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08896_ (.A1(_02476_),
    .A2(_03199_),
    .B(_03202_),
    .C(_02489_),
    .ZN(_03203_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08897_ (.A1(_02471_),
    .A2(_03196_),
    .B(_03203_),
    .C(_02518_),
    .ZN(_03204_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08898_ (.A1(_03195_),
    .A2(_03204_),
    .B(_02520_),
    .ZN(_03205_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08899_ (.A1(_02039_),
    .A2(_03186_),
    .A3(_03205_),
    .ZN(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08900_ (.I0(\mod.u_cpu.rf_ram.memory[512][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[513][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[514][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[515][1] ),
    .S0(_02494_),
    .S1(_02495_),
    .Z(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08901_ (.I(\mod.u_cpu.rf_ram.memory[517][1] ),
    .ZN(_03208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08902_ (.A1(_02507_),
    .A2(_03208_),
    .ZN(_03209_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08903_ (.A1(_02527_),
    .A2(\mod.u_cpu.rf_ram.memory[516][1] ),
    .B(_03209_),
    .ZN(_03210_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08904_ (.I(\mod.u_cpu.rf_ram.memory[519][1] ),
    .ZN(_03211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08905_ (.A1(_02500_),
    .A2(_03211_),
    .ZN(_03212_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08906_ (.A1(_02533_),
    .A2(\mod.u_cpu.rf_ram.memory[518][1] ),
    .B(_03212_),
    .C(_02537_),
    .ZN(_03213_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08907_ (.A1(_02525_),
    .A2(_03210_),
    .B(_03213_),
    .C(_02467_),
    .ZN(_03214_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08908_ (.A1(_02449_),
    .A2(_03207_),
    .B(_03214_),
    .C(_02469_),
    .ZN(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08909_ (.I0(\mod.u_cpu.rf_ram.memory[520][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[521][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[522][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[523][1] ),
    .S0(_02507_),
    .S1(_02543_),
    .Z(_03216_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08910_ (.I(\mod.u_cpu.rf_ram.memory[525][1] ),
    .ZN(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08911_ (.A1(_02509_),
    .A2(_03217_),
    .ZN(_03218_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08912_ (.A1(_02546_),
    .A2(\mod.u_cpu.rf_ram.memory[524][1] ),
    .B(_03218_),
    .ZN(_03219_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08913_ (.I(\mod.u_cpu.rf_ram.memory[527][1] ),
    .ZN(_03220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08914_ (.A1(_02551_),
    .A2(_03220_),
    .ZN(_03221_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08915_ (.A1(_02550_),
    .A2(\mod.u_cpu.rf_ram.memory[526][1] ),
    .B(_03221_),
    .C(_02515_),
    .ZN(_03222_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08916_ (.A1(_02545_),
    .A2(_03219_),
    .B(_03222_),
    .C(_02489_),
    .ZN(_03223_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08917_ (.A1(_02471_),
    .A2(_03216_),
    .B(_03223_),
    .C(_02491_),
    .ZN(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08918_ (.A1(_03215_),
    .A2(_03224_),
    .B(_01447_),
    .ZN(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08919_ (.I0(\mod.u_cpu.rf_ram.memory[536][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[537][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[538][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[539][1] ),
    .S0(_02560_),
    .S1(_02495_),
    .Z(_03226_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08920_ (.I(\mod.u_cpu.rf_ram.memory[541][1] ),
    .ZN(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08921_ (.A1(_02528_),
    .A2(_03227_),
    .ZN(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08922_ (.A1(_02527_),
    .A2(\mod.u_cpu.rf_ram.memory[540][1] ),
    .B(_03228_),
    .ZN(_03229_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08923_ (.I(\mod.u_cpu.rf_ram.memory[543][1] ),
    .ZN(_03230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08924_ (.A1(_02534_),
    .A2(_03230_),
    .ZN(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08925_ (.A1(_02533_),
    .A2(\mod.u_cpu.rf_ram.memory[542][1] ),
    .B(_03231_),
    .C(_02537_),
    .ZN(_03232_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08926_ (.A1(_02525_),
    .A2(_03229_),
    .B(_03232_),
    .C(_02539_),
    .ZN(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08927_ (.A1(_02523_),
    .A2(_03226_),
    .B(_03233_),
    .C(_02505_),
    .ZN(_03234_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08928_ (.I0(\mod.u_cpu.rf_ram.memory[528][1] ),
    .I1(\mod.u_cpu.rf_ram.memory[529][1] ),
    .I2(\mod.u_cpu.rf_ram.memory[530][1] ),
    .I3(\mod.u_cpu.rf_ram.memory[531][1] ),
    .S0(_02528_),
    .S1(_02543_),
    .Z(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08929_ (.I(\mod.u_cpu.rf_ram.memory[533][1] ),
    .ZN(_03236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08930_ (.A1(_02509_),
    .A2(_03236_),
    .ZN(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08931_ (.A1(_02546_),
    .A2(\mod.u_cpu.rf_ram.memory[532][1] ),
    .B(_03237_),
    .ZN(_03238_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08932_ (.I(\mod.u_cpu.rf_ram.memory[535][1] ),
    .ZN(_03239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08933_ (.A1(_02551_),
    .A2(_03239_),
    .ZN(_03240_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08934_ (.A1(_02550_),
    .A2(\mod.u_cpu.rf_ram.memory[534][1] ),
    .B(_03240_),
    .C(_02515_),
    .ZN(_03241_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08935_ (.A1(_02545_),
    .A2(_03238_),
    .B(_03241_),
    .C(_02555_),
    .ZN(_03242_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08936_ (.A1(_02542_),
    .A2(_03235_),
    .B(_03242_),
    .C(_02518_),
    .ZN(_03243_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08937_ (.A1(_03234_),
    .A2(_03243_),
    .B(_02520_),
    .ZN(_03244_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08938_ (.A1(_01459_),
    .A2(_03225_),
    .A3(_03244_),
    .ZN(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _08939_ (.A1(_01464_),
    .A2(_01465_),
    .A3(_03206_),
    .A4(_03245_),
    .Z(_03246_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _08940_ (.A1(_01466_),
    .A2(_02914_),
    .A3(_03167_),
    .B(_03246_),
    .ZN(_00001_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08941_ (.I(\mod.u_cpu.rf_ram.rdata[0] ),
    .ZN(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08942_ (.A1(_03247_),
    .A2(\mod.u_cpu.rf_ram.regzero ),
    .ZN(_03248_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08943_ (.I0(\mod.u_cpu.rf_ram_if.rdata0[1] ),
    .I1(_03248_),
    .S(_01478_),
    .Z(_03249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08944_ (.I(_03249_),
    .Z(_00002_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08945_ (.I(_01440_),
    .Z(_03250_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08946_ (.I(_01421_),
    .Z(_03251_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08947_ (.I(_03251_),
    .ZN(_03252_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08948_ (.I(_01422_),
    .Z(_03253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08949_ (.I(\mod.u_cpu.cpu.decode.opcode[0] ),
    .Z(_03254_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08950_ (.I(_03254_),
    .ZN(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08951_ (.A1(_03252_),
    .A2(_03253_),
    .A3(_03255_),
    .ZN(_03256_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08952_ (.I(_03256_),
    .ZN(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08953_ (.A1(\mod.u_cpu.cpu.mem_bytecnt[0] ),
    .A2(\mod.u_cpu.cpu.state.o_cnt[2] ),
    .A3(\mod.u_cpu.cpu.mem_bytecnt[1] ),
    .ZN(_03258_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08954_ (.I(_03258_),
    .Z(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08955_ (.A1(\mod.u_cpu.cpu.state.o_cnt_r[0] ),
    .A2(_03259_),
    .ZN(_03260_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08956_ (.I(\mod.u_arbiter.i_wb_cpu_dbus_we ),
    .Z(_03261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08957_ (.A1(\mod.u_cpu.cpu.decode.co_ebreak ),
    .A2(_01423_),
    .ZN(_03262_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08958_ (.A1(\mod.u_cpu.cpu.decode.opcode[2] ),
    .A2(\mod.u_cpu.cpu.decode.opcode[0] ),
    .A3(\mod.u_cpu.cpu.decode.opcode[1] ),
    .ZN(_03263_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08959_ (.A1(_03254_),
    .A2(\mod.u_cpu.cpu.decode.opcode[1] ),
    .B(_03263_),
    .ZN(_03264_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08960_ (.A1(_03253_),
    .A2(_03261_),
    .B(_03262_),
    .C(_03264_),
    .ZN(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08961_ (.A1(\mod.u_arbiter.i_wb_cpu_ibus_adr[0] ),
    .A2(_03265_),
    .ZN(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08962_ (.A1(\mod.u_cpu.cpu.ctrl.pc_plus_offset_cy_r ),
    .A2(_03266_),
    .Z(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08963_ (.I(\mod.u_cpu.cpu.mem_bytecnt[1] ),
    .Z(_03268_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08964_ (.I(\mod.u_cpu.cpu.mem_bytecnt[0] ),
    .Z(_03269_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08965_ (.A1(_03269_),
    .A2(\mod.u_cpu.cpu.state.o_cnt[2] ),
    .Z(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08966_ (.I(\mod.u_cpu.cpu.immdec.imm11_7[0] ),
    .ZN(_03271_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08967_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_we ),
    .A2(_03271_),
    .A3(_03263_),
    .Z(_03272_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08968_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_we ),
    .A2(_03263_),
    .B(\mod.u_cpu.cpu.immdec.imm24_20[0] ),
    .ZN(_03273_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08969_ (.A1(_01421_),
    .A2(\mod.u_cpu.cpu.branch_op ),
    .A3(\mod.u_cpu.cpu.csr_d_sel ),
    .ZN(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08970_ (.A1(\mod.u_cpu.cpu.bufreg2.i_cnt_done ),
    .A2(\mod.u_cpu.cpu.immdec.imm31 ),
    .A3(_03274_),
    .ZN(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _08971_ (.A1(\mod.u_cpu.cpu.bufreg2.i_cnt_done ),
    .A2(_03272_),
    .A3(_03273_),
    .B(_03275_),
    .ZN(_03276_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08972_ (.A1(_03268_),
    .A2(_03270_),
    .B(_03276_),
    .ZN(_03277_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08973_ (.A1(_03256_),
    .A2(_03277_),
    .Z(_03278_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08974_ (.I(\mod.u_cpu.cpu.bufreg.lsb[0] ),
    .Z(_03279_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08975_ (.I(\mod.u_cpu.cpu.decode.co_mem_word ),
    .ZN(_03280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08976_ (.A1(_03251_),
    .A2(_03280_),
    .ZN(_03281_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08977_ (.I(\mod.u_cpu.cpu.state.stage_two_req ),
    .ZN(_03282_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08978_ (.A1(_01430_),
    .A2(\mod.u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .B(\mod.u_cpu.cpu.state.init_done ),
    .C(_03282_),
    .ZN(_03283_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08979_ (.I(\mod.u_cpu.cpu.state.init_done ),
    .ZN(_03284_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _08980_ (.A1(\mod.u_cpu.cpu.state.genblk1.misalign_trap_sync_r ),
    .A2(_03284_),
    .A3(\mod.u_cpu.cpu.genblk3.csr.o_new_irq ),
    .A4(_01422_),
    .ZN(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08981_ (.A1(_01428_),
    .A2(_01429_),
    .ZN(_03286_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08982_ (.A1(\mod.u_cpu.cpu.decode.co_mem_word ),
    .A2(\mod.u_cpu.cpu.csr_d_sel ),
    .Z(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08983_ (.A1(\mod.u_cpu.cpu.branch_op ),
    .A2(_03254_),
    .Z(_03288_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _08984_ (.A1(_03286_),
    .A2(_03287_),
    .A3(_03288_),
    .B(_01421_),
    .ZN(_03289_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _08985_ (.A1(\mod.u_cpu.cpu.state.o_cnt_r[1] ),
    .A2(\mod.u_cpu.cpu.state.o_cnt_r[0] ),
    .A3(\mod.u_cpu.cpu.state.o_cnt_r[3] ),
    .A4(\mod.u_cpu.cpu.state.o_cnt_r[2] ),
    .Z(_03290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08986_ (.A1(_03289_),
    .A2(_03290_),
    .ZN(_03291_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _08987_ (.A1(_03281_),
    .A2(_03283_),
    .B1(_03285_),
    .B2(_03291_),
    .ZN(_03292_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08988_ (.A1(_03279_),
    .A2(_03292_),
    .B(_03256_),
    .ZN(_03293_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _08989_ (.A1(_03267_),
    .A2(_03278_),
    .A3(_03293_),
    .Z(_03294_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08990_ (.A1(_03278_),
    .A2(_03293_),
    .B(_03267_),
    .ZN(_03295_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08991_ (.A1(_03260_),
    .A2(_03294_),
    .A3(_03295_),
    .ZN(_03296_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08992_ (.I(_03251_),
    .Z(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08993_ (.I(_03253_),
    .ZN(_03298_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08994_ (.I(\mod.u_cpu.cpu.bne_or_bge ),
    .ZN(_03299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08995_ (.A1(_03280_),
    .A2(_03299_),
    .ZN(_03300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _08996_ (.A1(_03261_),
    .A2(\mod.u_cpu.cpu.bufreg.i_sh_signed ),
    .B(_03300_),
    .C(_01422_),
    .ZN(_03301_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08997_ (.I0(\mod.u_cpu.rf_ram_if.rdata1 ),
    .I1(_03248_),
    .S(\mod.u_cpu.rf_ram_if.rtrig1 ),
    .Z(_03302_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08998_ (.I0(_03276_),
    .I1(_03302_),
    .S(_03261_),
    .Z(_03303_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08999_ (.A1(_03301_),
    .A2(_03303_),
    .Z(_03304_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09000_ (.A1(\mod.u_cpu.cpu.alu.add_cy_r ),
    .A2(\mod.u_cpu.cpu.alu.i_rs1 ),
    .A3(_03304_),
    .Z(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09001_ (.I(_03299_),
    .Z(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09002_ (.I(_01430_),
    .Z(_03307_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09003_ (.I(\mod.u_cpu.cpu.alu.i_rs1 ),
    .Z(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09004_ (.I(_03303_),
    .Z(_03309_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09005_ (.A1(_03308_),
    .A2(_03309_),
    .Z(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09006_ (.A1(_03306_),
    .A2(_03307_),
    .A3(_03310_),
    .ZN(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09007_ (.A1(_03308_),
    .A2(_03309_),
    .Z(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09008_ (.I(\mod.u_cpu.cpu.alu.cmp_r ),
    .ZN(_03313_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09009_ (.A1(_01430_),
    .A2(_03313_),
    .A3(_03260_),
    .ZN(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09010_ (.I(_01428_),
    .Z(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09011_ (.A1(\mod.u_cpu.cpu.bufreg.lsb[0] ),
    .A2(_03292_),
    .Z(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09012_ (.A1(_03312_),
    .A2(_03287_),
    .B1(_03314_),
    .B2(_03315_),
    .C(_03316_),
    .ZN(_03317_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09013_ (.A1(_01431_),
    .A2(_03305_),
    .B(_03311_),
    .C(_03317_),
    .ZN(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09014_ (.A1(_03297_),
    .A2(_03298_),
    .A3(_03255_),
    .A4(_03318_),
    .ZN(_03319_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09015_ (.I(\mod.u_cpu.cpu.state.o_cnt_r[1] ),
    .ZN(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09016_ (.A1(\mod.u_cpu.cpu.state.o_cnt_r[2] ),
    .A2(\mod.u_cpu.cpu.ctrl.i_iscomp ),
    .ZN(_03321_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09017_ (.A1(_03320_),
    .A2(\mod.u_cpu.cpu.ctrl.i_iscomp ),
    .B(_03321_),
    .ZN(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09018_ (.A1(_03259_),
    .A2(_03322_),
    .Z(_03323_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09019_ (.A1(\mod.u_arbiter.i_wb_cpu_ibus_adr[0] ),
    .A2(\mod.u_cpu.cpu.ctrl.pc_plus_4_cy_r ),
    .Z(_03324_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09020_ (.A1(_03323_),
    .A2(_03324_),
    .Z(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09021_ (.A1(_03298_),
    .A2(_03255_),
    .ZN(_03326_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09022_ (.I(\mod.u_cpu.cpu.mem_if.signbit ),
    .ZN(_03327_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09023_ (.A1(_03306_),
    .A2(_03269_),
    .B(_03268_),
    .ZN(_03328_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _09024_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_dat[0] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_dat[16] ),
    .I2(\mod.u_arbiter.i_wb_cpu_dbus_dat[8] ),
    .I3(\mod.u_arbiter.i_wb_cpu_dbus_dat[24] ),
    .S0(\mod.u_cpu.cpu.bufreg.lsb[1] ),
    .S1(\mod.u_cpu.cpu.bufreg.lsb[0] ),
    .Z(_03329_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09025_ (.A1(_01428_),
    .A2(_03328_),
    .B(_03329_),
    .ZN(_03330_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09026_ (.A1(_03315_),
    .A2(_03327_),
    .A3(_03328_),
    .B(_03330_),
    .ZN(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09027_ (.I(_03254_),
    .Z(_03331_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09028_ (.A1(_03307_),
    .A2(_03330_),
    .B(_03251_),
    .C(_03331_),
    .ZN(_03332_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09029_ (.I(_03302_),
    .ZN(_03333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09030_ (.I(_03290_),
    .Z(_03334_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09031_ (.A1(_01435_),
    .A2(\mod.u_cpu.cpu.decode.co_ebreak ),
    .A3(_01452_),
    .ZN(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09032_ (.A1(_03334_),
    .A2(_03335_),
    .Z(_03336_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09033_ (.I(_03258_),
    .Z(_03337_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09034_ (.I(\mod.u_cpu.cpu.bufreg2.i_cnt_done ),
    .Z(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09035_ (.A1(_03338_),
    .A2(\mod.u_cpu.cpu.genblk3.csr.mcause31 ),
    .ZN(_03339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09036_ (.A1(\mod.u_cpu.cpu.genblk3.csr.mcause3_0[0] ),
    .A2(_03259_),
    .ZN(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09037_ (.A1(_03337_),
    .A2(_03339_),
    .B(_03340_),
    .ZN(_03341_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09038_ (.I(\mod.u_cpu.cpu.decode.op22 ),
    .ZN(_03342_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09039_ (.A1(\mod.u_cpu.cpu.decode.op26 ),
    .A2(_01452_),
    .ZN(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09040_ (.A1(\mod.u_cpu.cpu.state.o_cnt_r[3] ),
    .A2(_03342_),
    .A3(_03259_),
    .A4(_03343_),
    .Z(_03344_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09041_ (.A1(_03336_),
    .A2(_03341_),
    .B1(_03344_),
    .B2(\mod.u_cpu.cpu.genblk3.csr.mstatus_mie ),
    .ZN(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09042_ (.A1(_01432_),
    .A2(_03333_),
    .B(_03345_),
    .ZN(_03346_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09043_ (.A1(_03325_),
    .A2(_03326_),
    .B1(_01394_),
    .B2(_03332_),
    .C(_03346_),
    .ZN(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09044_ (.A1(_03257_),
    .A2(_03296_),
    .B(_03319_),
    .C(_03347_),
    .ZN(_03348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09045_ (.I(_03253_),
    .Z(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09046_ (.A1(_03349_),
    .A2(_03316_),
    .ZN(_03350_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09047_ (.A1(_03349_),
    .A2(_03296_),
    .B(_03350_),
    .C(_03250_),
    .ZN(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09048_ (.A1(_03250_),
    .A2(_03348_),
    .B(_03351_),
    .ZN(_03352_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09049_ (.I(_03352_),
    .ZN(\mod.u_cpu.cpu.o_wdata0 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09050_ (.I(_03250_),
    .Z(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09051_ (.I(_03307_),
    .Z(_03354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09052_ (.I(_03354_),
    .Z(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09053_ (.I(_03308_),
    .Z(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09054_ (.I(_03356_),
    .ZN(_03357_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09055_ (.A1(_03354_),
    .A2(_03357_),
    .ZN(_03358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09056_ (.I(_03280_),
    .Z(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09057_ (.A1(_03355_),
    .A2(\mod.u_cpu.cpu.csr_imm ),
    .B(_03358_),
    .C(_03359_),
    .ZN(_03360_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09058_ (.A1(_03306_),
    .A2(_03360_),
    .B(_03346_),
    .ZN(_03361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09059_ (.I(_03315_),
    .Z(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09060_ (.I(_01429_),
    .Z(_03363_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09061_ (.I(\mod.u_cpu.cpu.csr_imm ),
    .ZN(_03364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09062_ (.I(_03356_),
    .Z(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09063_ (.A1(_03354_),
    .A2(_03365_),
    .ZN(_03366_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09064_ (.A1(_03362_),
    .A2(_03363_),
    .B1(_03355_),
    .B2(_03364_),
    .C(_03366_),
    .ZN(_03367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09065_ (.A1(_03300_),
    .A2(_03367_),
    .ZN(_03368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09066_ (.A1(_03361_),
    .A2(_03368_),
    .ZN(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09067_ (.A1(_03353_),
    .A2(_03369_),
    .ZN(_03370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09068_ (.I(\mod.u_arbiter.i_wb_cpu_ibus_adr[0] ),
    .Z(_03371_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09069_ (.I(_01433_),
    .ZN(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09070_ (.A1(_01434_),
    .A2(_01436_),
    .ZN(_03373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09071_ (.A1(_03372_),
    .A2(_03373_),
    .ZN(_03374_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09072_ (.I(_03374_),
    .Z(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09073_ (.A1(_03371_),
    .A2(_03375_),
    .ZN(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09074_ (.A1(_03370_),
    .A2(_03376_),
    .ZN(\mod.u_cpu.cpu.o_wdata1 ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09075_ (.I(_03334_),
    .Z(_03377_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09076_ (.I(_03377_),
    .Z(_03378_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09077_ (.A1(\mod.u_cpu.cpu.alu.add_cy_r ),
    .A2(_03308_),
    .ZN(_03379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09078_ (.A1(\mod.u_cpu.cpu.alu.add_cy_r ),
    .A2(_03356_),
    .ZN(_03380_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09079_ (.A1(_03379_),
    .A2(_03304_),
    .B(_03380_),
    .ZN(_03381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09080_ (.A1(_03378_),
    .A2(_03381_),
    .ZN(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09081_ (.A1(_03301_),
    .A2(_03378_),
    .B(_03382_),
    .ZN(_00003_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09082_ (.I(net1),
    .ZN(_03383_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09083_ (.I(net2),
    .ZN(_03384_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09084_ (.I(_03384_),
    .Z(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09085_ (.I(_03385_),
    .Z(_03386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09086_ (.I(_03386_),
    .Z(_03387_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09087_ (.I(\mod.u_cpu.cpu.state.o_cnt_r[0] ),
    .Z(_03388_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09088_ (.I(\mod.u_cpu.cpu.state.o_cnt_r[3] ),
    .Z(_03389_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09089_ (.A1(\mod.u_cpu.cpu.state.o_cnt_r[1] ),
    .A2(_03388_),
    .A3(_03389_),
    .A4(\mod.u_cpu.cpu.state.o_cnt_r[2] ),
    .ZN(_03390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09090_ (.I(_03390_),
    .Z(_03391_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09091_ (.I(\mod.u_cpu.cpu.bufreg.lsb[1] ),
    .Z(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09092_ (.A1(_03362_),
    .A2(_03392_),
    .B1(_03300_),
    .B2(_03279_),
    .ZN(_03393_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09093_ (.I(_03297_),
    .Z(_03394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09094_ (.I(_03349_),
    .Z(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09095_ (.A1(_03394_),
    .A2(_03395_),
    .ZN(_03396_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09096_ (.A1(\mod.u_cpu.cpu.state.init_done ),
    .A2(_03391_),
    .A3(_03393_),
    .A4(_03396_),
    .ZN(_03397_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09097_ (.I(net5),
    .ZN(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09098_ (.A1(_03398_),
    .A2(\mod.u_cpu.cpu.state.ibus_cyc ),
    .Z(_03399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09099_ (.I(_03399_),
    .Z(_03400_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09100_ (.A1(_03385_),
    .A2(_03400_),
    .ZN(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09101_ (.I(_03401_),
    .Z(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09102_ (.A1(_03383_),
    .A2(_03387_),
    .B1(_03397_),
    .B2(_03402_),
    .ZN(_00008_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09103_ (.I(_03261_),
    .Z(_03403_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09104_ (.I(_03403_),
    .ZN(_03404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09105_ (.I(net2),
    .Z(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09106_ (.A1(_03398_),
    .A2(\mod.u_cpu.cpu.state.ibus_cyc ),
    .ZN(_03406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09107_ (.A1(_03405_),
    .A2(_03406_),
    .ZN(_03407_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09108_ (.I(_03407_),
    .Z(_03408_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09109_ (.I(_03385_),
    .Z(_03409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09110_ (.I(_03409_),
    .Z(_03410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09111_ (.A1(_03410_),
    .A2(\mod.timer_irq ),
    .ZN(_03411_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09112_ (.A1(_03404_),
    .A2(_03408_),
    .B(_03411_),
    .ZN(_00019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09113_ (.I(\mod.u_arbiter.i_wb_cpu_ack ),
    .Z(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09114_ (.I(_03405_),
    .Z(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09115_ (.I(_03413_),
    .Z(_03414_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09116_ (.I(_03414_),
    .Z(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09117_ (.I(_03279_),
    .Z(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09118_ (.I(_03413_),
    .Z(_03417_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09119_ (.A1(_03416_),
    .A2(_03392_),
    .B(_03417_),
    .ZN(_03418_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09120_ (.A1(_03412_),
    .A2(_03415_),
    .B(_03418_),
    .ZN(_03419_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09121_ (.I(_03419_),
    .ZN(_00030_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09122_ (.A1(_03363_),
    .A2(_03416_),
    .ZN(_03420_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09123_ (.A1(_03362_),
    .A2(_03385_),
    .ZN(_03421_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09124_ (.A1(_03392_),
    .A2(_03420_),
    .B(_03421_),
    .ZN(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09125_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[0] ),
    .A2(_03415_),
    .B(_03422_),
    .ZN(_03423_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09126_ (.I(_03423_),
    .ZN(_00041_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _09127_ (.I(\mod.u_arbiter.i_wb_cpu_rdt[1] ),
    .ZN(_03424_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09128_ (.I(_03416_),
    .ZN(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09129_ (.I(_03392_),
    .Z(_03426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09130_ (.A1(_03425_),
    .A2(_03426_),
    .ZN(_03427_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09131_ (.A1(_03424_),
    .A2(_03387_),
    .B1(_03427_),
    .B2(_03421_),
    .ZN(_00052_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _09132_ (.I(\mod.u_arbiter.i_wb_cpu_rdt[2] ),
    .ZN(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09133_ (.A1(_03363_),
    .A2(_03416_),
    .B(_03426_),
    .ZN(_03429_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09134_ (.A1(_03428_),
    .A2(_03387_),
    .B1(_03421_),
    .B2(_03429_),
    .ZN(_00063_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09135_ (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[0] ),
    .Z(_03430_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09136_ (.I(_03430_),
    .ZN(_03431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09137_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[3] ),
    .A2(_03410_),
    .ZN(_03432_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09138_ (.A1(_03431_),
    .A2(_03387_),
    .B(_03432_),
    .ZN(_00074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09139_ (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[1] ),
    .Z(_03433_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09140_ (.I(_03433_),
    .ZN(_03434_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09141_ (.I(_03409_),
    .Z(_03435_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09142_ (.I(_03409_),
    .Z(_03436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09143_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[4] ),
    .A2(_03436_),
    .ZN(_03437_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09144_ (.A1(_03434_),
    .A2(_03435_),
    .B(_03437_),
    .ZN(_00075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09145_ (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[2] ),
    .Z(_03438_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09146_ (.I(_03405_),
    .Z(_03439_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09147_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[5] ),
    .I1(_03438_),
    .S(_03439_),
    .Z(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09148_ (.I(_03440_),
    .Z(_00076_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09149_ (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[3] ),
    .Z(_03441_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09150_ (.I(_03417_),
    .Z(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09151_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[6] ),
    .I1(_03441_),
    .S(_03442_),
    .Z(_03443_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09152_ (.I(_03443_),
    .Z(_00077_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09153_ (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[4] ),
    .Z(_03444_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09154_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[7] ),
    .I1(_03444_),
    .S(_03442_),
    .Z(_03445_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09155_ (.I(_03445_),
    .Z(_00009_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09156_ (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .ZN(_03446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09157_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[8] ),
    .A2(_03436_),
    .ZN(_03447_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09158_ (.A1(_03446_),
    .A2(_03435_),
    .B(_03447_),
    .ZN(_00010_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09159_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[9] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_dat[6] ),
    .S(_03442_),
    .Z(_03448_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09160_ (.I(_03448_),
    .Z(_00011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09161_ (.I(\mod.u_arbiter.i_wb_cpu_rdt[10] ),
    .Z(_03449_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09162_ (.I0(_03449_),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_dat[7] ),
    .S(_03442_),
    .Z(_03450_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09163_ (.I(_03450_),
    .Z(_00012_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09164_ (.I(_03413_),
    .Z(_03451_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09165_ (.I(_03451_),
    .Z(_03452_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09166_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[11] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_dat[8] ),
    .S(_03452_),
    .Z(_03453_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09167_ (.I(_03453_),
    .Z(_00013_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09168_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[12] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_dat[9] ),
    .S(_03452_),
    .Z(_03454_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09169_ (.I(_03454_),
    .Z(_00014_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09170_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[13] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_dat[10] ),
    .S(_03452_),
    .Z(_03455_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09171_ (.I(_03455_),
    .Z(_00015_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09172_ (.I(\mod.u_arbiter.i_wb_cpu_rdt[14] ),
    .Z(_03456_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09173_ (.I0(_03456_),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_dat[11] ),
    .S(_03452_),
    .Z(_03457_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09174_ (.I(_03457_),
    .Z(_00016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09175_ (.I(\mod.u_arbiter.i_wb_cpu_rdt[15] ),
    .Z(_03458_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09176_ (.I(_03451_),
    .Z(_03459_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09177_ (.I0(_03458_),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_dat[12] ),
    .S(_03459_),
    .Z(_03460_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09178_ (.I(_03460_),
    .Z(_00017_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09179_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[16] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_dat[13] ),
    .S(_03459_),
    .Z(_03461_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09180_ (.I(_03461_),
    .Z(_00018_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09181_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[17] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_dat[14] ),
    .S(_03459_),
    .Z(_03462_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09182_ (.I(_03462_),
    .Z(_00020_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09183_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[18] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_dat[15] ),
    .S(_03459_),
    .Z(_03463_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09184_ (.I(_03463_),
    .Z(_00021_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09185_ (.I(_03451_),
    .Z(_03464_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09186_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[19] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_dat[16] ),
    .S(_03464_),
    .Z(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09187_ (.I(_03465_),
    .Z(_00022_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09188_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[20] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_dat[17] ),
    .S(_03464_),
    .Z(_03466_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09189_ (.I(_03466_),
    .Z(_00023_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09190_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[21] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_dat[18] ),
    .S(_03464_),
    .Z(_03467_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09191_ (.I(_03467_),
    .Z(_00024_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09192_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[22] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_dat[19] ),
    .S(_03464_),
    .Z(_03468_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09193_ (.I(_03468_),
    .Z(_00025_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09194_ (.I(_03451_),
    .Z(_03469_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09195_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[23] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_dat[20] ),
    .S(_03469_),
    .Z(_03470_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09196_ (.I(_03470_),
    .Z(_00026_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09197_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[24] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_dat[21] ),
    .S(_03469_),
    .Z(_03471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09198_ (.I(_03471_),
    .Z(_00027_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09199_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[25] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_dat[22] ),
    .S(_03469_),
    .Z(_03472_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09200_ (.I(_03472_),
    .Z(_00028_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09201_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[26] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_dat[23] ),
    .S(_03469_),
    .Z(_03473_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09202_ (.I(_03473_),
    .Z(_00029_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09203_ (.I(_03414_),
    .Z(_03474_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09204_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[27] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_dat[24] ),
    .S(_03474_),
    .Z(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09205_ (.I(_03475_),
    .Z(_00031_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09206_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[28] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_dat[25] ),
    .S(_03474_),
    .Z(_03476_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09207_ (.I(_03476_),
    .Z(_00032_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09208_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[29] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_dat[26] ),
    .S(_03474_),
    .Z(_03477_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09209_ (.I(_03477_),
    .Z(_00033_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09210_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[30] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_dat[27] ),
    .S(_03474_),
    .Z(_03478_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09211_ (.I(_03478_),
    .Z(_00034_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09212_ (.I(_03414_),
    .Z(_03479_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09213_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[31] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_dat[28] ),
    .S(_03479_),
    .Z(_03480_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09214_ (.I(_03480_),
    .Z(_00035_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09215_ (.I0(\mod.u_scanchain_local.module_data_in[34] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_dat[29] ),
    .S(_03479_),
    .Z(_03481_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09216_ (.I(_03481_),
    .Z(_00036_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09217_ (.I0(\mod.u_scanchain_local.module_data_in[35] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_dat[30] ),
    .S(_03479_),
    .Z(_03482_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09218_ (.I(_03482_),
    .Z(_00037_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09219_ (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[31] ),
    .ZN(_03483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09220_ (.A1(_03410_),
    .A2(\mod.u_scanchain_local.module_data_in[36] ),
    .ZN(_03484_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09221_ (.A1(_03483_),
    .A2(_03435_),
    .B(_03484_),
    .ZN(_00038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09222_ (.A1(_03435_),
    .A2(\mod.u_scanchain_local.module_data_in[37] ),
    .ZN(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09223_ (.I(_03406_),
    .Z(_03486_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09224_ (.A1(_03384_),
    .A2(_03486_),
    .ZN(_03487_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09225_ (.I(_03487_),
    .Z(_03488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09226_ (.I(_03488_),
    .Z(_03489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09227_ (.A1(_03371_),
    .A2(_03489_),
    .ZN(_03490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09228_ (.A1(_03485_),
    .A2(_03490_),
    .ZN(_00039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09229_ (.A1(_03410_),
    .A2(\mod.u_scanchain_local.module_data_in[38] ),
    .ZN(_03491_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09230_ (.I(\mod.u_arbiter.i_wb_cpu_ibus_adr[1] ),
    .Z(_03492_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09231_ (.I(_03487_),
    .Z(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09232_ (.A1(_03492_),
    .A2(_03493_),
    .ZN(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09233_ (.A1(_03491_),
    .A2(_03494_),
    .ZN(_00040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09234_ (.I(_03405_),
    .Z(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09235_ (.I(_03495_),
    .Z(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09236_ (.A1(_03414_),
    .A2(_03400_),
    .ZN(_03497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09237_ (.I(\mod.u_cpu.cpu.genblk1.align.ctrl_misal ),
    .Z(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09238_ (.I(_03498_),
    .Z(_03499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09239_ (.I(_03499_),
    .Z(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09240_ (.I(_03500_),
    .Z(_03501_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09241_ (.I(_03501_),
    .Z(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09242_ (.I(_03502_),
    .Z(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09243_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[2] ),
    .A2(_03503_),
    .Z(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _09244_ (.A1(_03496_),
    .A2(\mod.u_scanchain_local.module_data_in[39] ),
    .B1(_03497_),
    .B2(_03504_),
    .C1(_03408_),
    .C2(\mod.u_arbiter.i_wb_cpu_dbus_adr[2] ),
    .ZN(_03505_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09245_ (.I(_03505_),
    .ZN(_00042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09246_ (.I(_03493_),
    .Z(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09247_ (.I(\mod.u_cpu.cpu.ctrl.o_ibus_adr[3] ),
    .Z(_03507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09248_ (.I(\mod.u_cpu.cpu.ctrl.o_ibus_adr[2] ),
    .Z(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09249_ (.I(_03502_),
    .Z(_03509_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09250_ (.I(_03509_),
    .Z(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09251_ (.A1(_03508_),
    .A2(_03510_),
    .ZN(_03511_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09252_ (.A1(_03507_),
    .A2(_03511_),
    .Z(_03512_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09253_ (.A1(_03479_),
    .A2(\mod.u_scanchain_local.module_data_in[40] ),
    .B1(_03408_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_adr[3] ),
    .ZN(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09254_ (.A1(_03506_),
    .A2(_03512_),
    .B(_03513_),
    .ZN(_00043_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09255_ (.A1(_03507_),
    .A2(_03508_),
    .A3(_03503_),
    .ZN(_03514_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09256_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[4] ),
    .A2(_03514_),
    .Z(_03515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09257_ (.I(_03495_),
    .Z(_03516_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09258_ (.I(_03407_),
    .Z(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09259_ (.I(_03517_),
    .Z(_03518_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09260_ (.A1(_03516_),
    .A2(\mod.u_scanchain_local.module_data_in[41] ),
    .B1(_03518_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_adr[4] ),
    .ZN(_03519_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09261_ (.A1(_03506_),
    .A2(_03515_),
    .B(_03519_),
    .ZN(_00044_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09262_ (.I(\mod.u_cpu.cpu.ctrl.o_ibus_adr[5] ),
    .Z(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09263_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[4] ),
    .A2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[3] ),
    .A3(\mod.u_cpu.cpu.ctrl.o_ibus_adr[2] ),
    .A4(_03498_),
    .Z(_03521_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09264_ (.A1(_03520_),
    .A2(_03521_),
    .ZN(_03522_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09265_ (.A1(_03516_),
    .A2(\mod.u_scanchain_local.module_data_in[42] ),
    .B1(_03518_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_adr[5] ),
    .ZN(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09266_ (.A1(_03506_),
    .A2(_03522_),
    .B(_03523_),
    .ZN(_00045_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09267_ (.I(\mod.u_cpu.cpu.ctrl.o_ibus_adr[6] ),
    .Z(_03524_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09268_ (.A1(_03520_),
    .A2(_03521_),
    .Z(_03525_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09269_ (.A1(_03524_),
    .A2(_03525_),
    .ZN(_03526_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09270_ (.A1(_03516_),
    .A2(\mod.u_scanchain_local.module_data_in[43] ),
    .B1(_03518_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_adr[6] ),
    .ZN(_03527_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09271_ (.A1(_03506_),
    .A2(_03526_),
    .B(_03527_),
    .ZN(_00046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09272_ (.I(_03488_),
    .Z(_03528_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09273_ (.A1(_03524_),
    .A2(_03525_),
    .ZN(_03529_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09274_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[7] ),
    .A2(_03529_),
    .Z(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09275_ (.A1(_03516_),
    .A2(\mod.u_scanchain_local.module_data_in[44] ),
    .B1(_03518_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_adr[7] ),
    .ZN(_03531_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09276_ (.A1(_03528_),
    .A2(_03530_),
    .B(_03531_),
    .ZN(_00047_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09277_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[7] ),
    .A2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[6] ),
    .Z(_03532_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09278_ (.A1(_03525_),
    .A2(_03532_),
    .ZN(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09279_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[8] ),
    .A2(_03533_),
    .Z(_03534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09280_ (.I(_03495_),
    .Z(_03535_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09281_ (.I(_03517_),
    .Z(_03536_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09282_ (.A1(_03535_),
    .A2(\mod.u_scanchain_local.module_data_in[45] ),
    .B1(_03536_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_adr[8] ),
    .ZN(_03537_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09283_ (.A1(_03528_),
    .A2(_03534_),
    .B(_03537_),
    .ZN(_00048_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _09284_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[8] ),
    .A2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[5] ),
    .A3(_03521_),
    .A4(_03532_),
    .ZN(_03538_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09285_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[9] ),
    .A2(_03538_),
    .Z(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09286_ (.A1(_03535_),
    .A2(\mod.u_scanchain_local.module_data_in[46] ),
    .B1(_03536_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_adr[9] ),
    .ZN(_03540_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09287_ (.A1(_03528_),
    .A2(_03539_),
    .B(_03540_),
    .ZN(_00049_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09288_ (.I(\mod.u_cpu.cpu.ctrl.o_ibus_adr[10] ),
    .Z(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _09289_ (.I(\mod.u_cpu.cpu.ctrl.o_ibus_adr[9] ),
    .ZN(_03542_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09290_ (.A1(_03542_),
    .A2(_03538_),
    .ZN(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09291_ (.A1(_03541_),
    .A2(_03543_),
    .ZN(_03544_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09292_ (.A1(_03535_),
    .A2(\mod.u_scanchain_local.module_data_in[47] ),
    .B1(_03536_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_adr[10] ),
    .ZN(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09293_ (.A1(_03528_),
    .A2(_03544_),
    .B(_03545_),
    .ZN(_00050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09294_ (.I(_03488_),
    .Z(_03546_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09295_ (.I(\mod.u_cpu.cpu.ctrl.o_ibus_adr[11] ),
    .Z(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09296_ (.A1(_03541_),
    .A2(_03543_),
    .Z(_03548_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09297_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[11] ),
    .A2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[10] ),
    .A3(_03543_),
    .ZN(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09298_ (.A1(_03547_),
    .A2(_03548_),
    .B(_03549_),
    .ZN(_03550_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09299_ (.A1(_03535_),
    .A2(\mod.u_scanchain_local.module_data_in[48] ),
    .B1(_03536_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_adr[11] ),
    .ZN(_03551_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09300_ (.A1(_03546_),
    .A2(_03550_),
    .B(_03551_),
    .ZN(_00051_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09301_ (.I(\mod.u_cpu.cpu.ctrl.o_ibus_adr[12] ),
    .Z(_03552_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09302_ (.A1(_03552_),
    .A2(_03549_),
    .Z(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09303_ (.I(_03495_),
    .Z(_03554_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09304_ (.I(_03407_),
    .Z(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09305_ (.A1(_03554_),
    .A2(\mod.u_scanchain_local.module_data_in[49] ),
    .B1(_03555_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_adr[12] ),
    .ZN(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09306_ (.A1(_03546_),
    .A2(_03553_),
    .B(_03556_),
    .ZN(_00053_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09307_ (.I(\mod.u_cpu.cpu.ctrl.o_ibus_adr[13] ),
    .ZN(_03557_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09308_ (.A1(_03552_),
    .A2(_03547_),
    .A3(\mod.u_cpu.cpu.ctrl.o_ibus_adr[10] ),
    .A4(_03543_),
    .ZN(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09309_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[13] ),
    .A2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[12] ),
    .ZN(_03559_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09310_ (.A1(_03549_),
    .A2(_03559_),
    .ZN(_03560_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09311_ (.I(_03486_),
    .Z(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09312_ (.A1(_03557_),
    .A2(_03558_),
    .B(_03560_),
    .C(_03561_),
    .ZN(_03562_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09313_ (.I(_03413_),
    .Z(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09314_ (.I(_03486_),
    .Z(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09315_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_adr[13] ),
    .A2(_03564_),
    .ZN(_03565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09316_ (.A1(_03563_),
    .A2(_03565_),
    .ZN(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09317_ (.A1(_03415_),
    .A2(\mod.u_scanchain_local.module_data_in[50] ),
    .B1(_03562_),
    .B2(_03566_),
    .ZN(_03567_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09318_ (.I(_03567_),
    .ZN(_00054_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09319_ (.I(_03497_),
    .Z(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09320_ (.I(\mod.u_cpu.cpu.ctrl.o_ibus_adr[14] ),
    .Z(_03569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09321_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[11] ),
    .A2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[10] ),
    .ZN(_03570_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _09322_ (.A1(_03542_),
    .A2(_03538_),
    .A3(_03570_),
    .A4(_03559_),
    .Z(_03571_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09323_ (.A1(_03569_),
    .A2(_03571_),
    .Z(_03572_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09324_ (.A1(_03436_),
    .A2(\mod.u_scanchain_local.module_data_in[51] ),
    .B1(_03402_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_adr[14] ),
    .ZN(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09325_ (.A1(_03568_),
    .A2(_03572_),
    .B(_03573_),
    .ZN(_00055_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09326_ (.I(\mod.u_cpu.cpu.ctrl.o_ibus_adr[15] ),
    .Z(_03574_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09327_ (.A1(_03569_),
    .A2(_03560_),
    .ZN(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09328_ (.A1(_03574_),
    .A2(_03575_),
    .Z(_03576_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09329_ (.A1(_03554_),
    .A2(\mod.u_scanchain_local.module_data_in[52] ),
    .B1(_03555_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_adr[15] ),
    .ZN(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09330_ (.A1(_03546_),
    .A2(_03576_),
    .B(_03577_),
    .ZN(_00056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09331_ (.I(\mod.u_cpu.cpu.ctrl.o_ibus_adr[16] ),
    .Z(_03578_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09332_ (.A1(_03574_),
    .A2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[14] ),
    .A3(_03560_),
    .ZN(_03579_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09333_ (.A1(_03578_),
    .A2(_03579_),
    .Z(_03580_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09334_ (.A1(_03554_),
    .A2(\mod.u_scanchain_local.module_data_in[53] ),
    .B1(_03555_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_adr[16] ),
    .ZN(_03581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09335_ (.A1(_03546_),
    .A2(_03580_),
    .B(_03581_),
    .ZN(_00057_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09336_ (.I(_03578_),
    .ZN(_03582_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09337_ (.A1(_03582_),
    .A2(_03579_),
    .ZN(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09338_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[17] ),
    .A2(_03583_),
    .ZN(_03584_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _09339_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[17] ),
    .A2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[16] ),
    .A3(\mod.u_cpu.cpu.ctrl.o_ibus_adr[15] ),
    .A4(\mod.u_cpu.cpu.ctrl.o_ibus_adr[14] ),
    .ZN(_03585_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09340_ (.A1(_03571_),
    .A2(_03585_),
    .ZN(_03586_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09341_ (.A1(_03386_),
    .A2(\mod.u_scanchain_local.module_data_in[54] ),
    .B1(_03401_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_adr[17] ),
    .ZN(_03587_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09342_ (.A1(_03568_),
    .A2(_03584_),
    .A3(_03586_),
    .B(_03587_),
    .ZN(_00058_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09343_ (.I(\mod.u_cpu.cpu.ctrl.o_ibus_adr[18] ),
    .Z(_03588_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09344_ (.A1(_03570_),
    .A2(_03559_),
    .Z(_03589_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09345_ (.A1(_03542_),
    .A2(_03538_),
    .A3(_03589_),
    .A4(_03585_),
    .ZN(_03590_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09346_ (.A1(_03588_),
    .A2(_03590_),
    .ZN(_03591_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09347_ (.A1(_03436_),
    .A2(\mod.u_scanchain_local.module_data_in[55] ),
    .B1(_03402_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_adr[18] ),
    .ZN(_03592_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09348_ (.A1(_03568_),
    .A2(_03591_),
    .B(_03592_),
    .ZN(_00059_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09349_ (.A1(_03588_),
    .A2(_03590_),
    .B(\mod.u_cpu.cpu.ctrl.o_ibus_adr[19] ),
    .ZN(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09350_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[19] ),
    .A2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[18] ),
    .Z(_03594_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09351_ (.A1(_03590_),
    .A2(_03594_),
    .Z(_03595_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09352_ (.A1(_03593_),
    .A2(_03595_),
    .B(_03488_),
    .ZN(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _09353_ (.A1(_03415_),
    .A2(\mod.u_scanchain_local.module_data_in[56] ),
    .B1(_03408_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_adr[19] ),
    .C(_03596_),
    .ZN(_03597_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09354_ (.I(_03597_),
    .ZN(_00060_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09355_ (.I(\mod.u_cpu.cpu.ctrl.o_ibus_adr[20] ),
    .Z(_03598_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09356_ (.A1(_03598_),
    .A2(_03586_),
    .A3(_03594_),
    .ZN(_03599_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09357_ (.A1(_03598_),
    .A2(_03595_),
    .B(_03599_),
    .ZN(_03600_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09358_ (.A1(_03554_),
    .A2(\mod.u_scanchain_local.module_data_in[57] ),
    .B1(_03555_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_adr[20] ),
    .ZN(_03601_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09359_ (.A1(_03489_),
    .A2(_03600_),
    .B(_03601_),
    .ZN(_00061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09360_ (.I(\mod.u_cpu.cpu.ctrl.o_ibus_adr[21] ),
    .Z(_03602_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09361_ (.A1(_03602_),
    .A2(_03599_),
    .Z(_03603_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09362_ (.A1(_03563_),
    .A2(\mod.u_scanchain_local.module_data_in[58] ),
    .B1(_03517_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_adr[21] ),
    .ZN(_03604_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09363_ (.A1(_03489_),
    .A2(_03603_),
    .B(_03604_),
    .ZN(_00062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09364_ (.I(\mod.u_cpu.cpu.ctrl.o_ibus_adr[22] ),
    .Z(_03605_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09365_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[21] ),
    .A2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[20] ),
    .A3(_03595_),
    .Z(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09366_ (.A1(_03605_),
    .A2(_03606_),
    .ZN(_03607_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09367_ (.A1(_03605_),
    .A2(_03606_),
    .Z(_03608_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09368_ (.A1(_03386_),
    .A2(\mod.u_scanchain_local.module_data_in[59] ),
    .B1(_03401_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_adr[22] ),
    .ZN(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09369_ (.A1(_03568_),
    .A2(_03607_),
    .A3(_03608_),
    .B(_03609_),
    .ZN(_00064_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09370_ (.I(\mod.u_cpu.cpu.ctrl.o_ibus_adr[23] ),
    .Z(_03610_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09371_ (.A1(_03610_),
    .A2(_03608_),
    .ZN(_03611_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09372_ (.A1(_03563_),
    .A2(\mod.u_scanchain_local.module_data_in[60] ),
    .B1(_03517_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_adr[23] ),
    .ZN(_03612_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09373_ (.A1(_03489_),
    .A2(_03611_),
    .B(_03612_),
    .ZN(_00065_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09374_ (.A1(_03496_),
    .A2(\mod.u_scanchain_local.module_data_in[61] ),
    .ZN(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09375_ (.I(_03486_),
    .Z(_03614_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09376_ (.I(_03614_),
    .Z(_03615_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09377_ (.I(\mod.u_cpu.cpu.ctrl.o_ibus_adr[24] ),
    .Z(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09378_ (.A1(_03610_),
    .A2(_03608_),
    .B(_03616_),
    .ZN(_03617_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09379_ (.A1(_03602_),
    .A2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[20] ),
    .A3(_03586_),
    .A4(_03594_),
    .ZN(_03618_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09380_ (.A1(_03616_),
    .A2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[23] ),
    .A3(\mod.u_cpu.cpu.ctrl.o_ibus_adr[22] ),
    .ZN(_03619_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09381_ (.A1(_03618_),
    .A2(_03619_),
    .ZN(_03620_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09382_ (.A1(_03564_),
    .A2(_03617_),
    .A3(_03620_),
    .B(_03417_),
    .ZN(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09383_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_adr[24] ),
    .A2(_03615_),
    .B(_03621_),
    .ZN(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09384_ (.A1(_03613_),
    .A2(_03622_),
    .ZN(_00066_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09385_ (.I(_03563_),
    .Z(_03623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09386_ (.I(\mod.u_cpu.cpu.ctrl.o_ibus_adr[25] ),
    .Z(_03624_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09387_ (.A1(_03624_),
    .A2(_03620_),
    .ZN(_03625_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09388_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[24] ),
    .A2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[23] ),
    .A3(\mod.u_cpu.cpu.ctrl.o_ibus_adr[22] ),
    .A4(_03606_),
    .Z(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09389_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[25] ),
    .A2(_03626_),
    .Z(_03627_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09390_ (.A1(_03564_),
    .A2(_03625_),
    .A3(_03627_),
    .ZN(_03628_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09391_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_adr[25] ),
    .A2(_03615_),
    .B(_03628_),
    .ZN(_03629_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09392_ (.A1(_03496_),
    .A2(\mod.u_scanchain_local.module_data_in[62] ),
    .ZN(_03630_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09393_ (.A1(_03623_),
    .A2(_03629_),
    .B(_03630_),
    .ZN(_00067_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09394_ (.I(\mod.u_cpu.cpu.ctrl.o_ibus_adr[26] ),
    .Z(_03631_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09395_ (.A1(_03631_),
    .A2(_03624_),
    .A3(_03620_),
    .Z(_03632_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09396_ (.A1(_03631_),
    .A2(_03627_),
    .B(_03493_),
    .ZN(_03633_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09397_ (.A1(_03386_),
    .A2(\mod.u_scanchain_local.module_data_in[63] ),
    .B1(_03401_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_adr[26] ),
    .ZN(_03634_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09398_ (.A1(_03632_),
    .A2(_03633_),
    .B(_03634_),
    .ZN(_00068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09399_ (.I(\mod.u_cpu.cpu.ctrl.o_ibus_adr[27] ),
    .Z(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09400_ (.A1(_03635_),
    .A2(_03632_),
    .ZN(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09401_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[27] ),
    .A2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[26] ),
    .A3(_03627_),
    .Z(_03637_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09402_ (.I(_03637_),
    .Z(_03638_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09403_ (.A1(_03614_),
    .A2(_03636_),
    .A3(_03638_),
    .ZN(_03639_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09404_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_adr[27] ),
    .A2(_03615_),
    .B(_03639_),
    .ZN(_03640_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09405_ (.A1(_03439_),
    .A2(\mod.u_scanchain_local.module_data_in[64] ),
    .ZN(_03641_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09406_ (.A1(_03623_),
    .A2(_03640_),
    .B(_03641_),
    .ZN(_00069_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09407_ (.I(\mod.u_cpu.cpu.ctrl.o_ibus_adr[28] ),
    .Z(_03642_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09408_ (.A1(_03642_),
    .A2(_03638_),
    .ZN(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09409_ (.A1(_03561_),
    .A2(_03643_),
    .ZN(_03644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09410_ (.A1(_03642_),
    .A2(_03638_),
    .ZN(_03645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09411_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_adr[28] ),
    .A2(_03561_),
    .B1(_03644_),
    .B2(_03645_),
    .ZN(_03646_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09412_ (.A1(_03439_),
    .A2(\mod.u_scanchain_local.module_data_in[65] ),
    .ZN(_03647_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09413_ (.A1(_03623_),
    .A2(_03646_),
    .B(_03647_),
    .ZN(_00070_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09414_ (.I(\mod.u_cpu.cpu.ctrl.o_ibus_adr[29] ),
    .Z(_03648_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09415_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[28] ),
    .A2(_03638_),
    .B(_03648_),
    .ZN(_03649_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09416_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[29] ),
    .A2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[28] ),
    .A3(_03635_),
    .A4(_03632_),
    .Z(_03650_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09417_ (.A1(_03614_),
    .A2(_03649_),
    .A3(_03650_),
    .ZN(_03651_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09418_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_adr[29] ),
    .A2(_03615_),
    .B(_03651_),
    .ZN(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09419_ (.A1(_03439_),
    .A2(\mod.u_scanchain_local.module_data_in[66] ),
    .ZN(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09420_ (.A1(_03623_),
    .A2(_03652_),
    .B(_03653_),
    .ZN(_00071_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09421_ (.A1(_03496_),
    .A2(\mod.u_scanchain_local.module_data_in[67] ),
    .ZN(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09422_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[30] ),
    .A2(_03650_),
    .ZN(_03655_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09423_ (.A1(_03564_),
    .A2(_03655_),
    .ZN(_03656_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09424_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[30] ),
    .A2(_03648_),
    .A3(\mod.u_cpu.cpu.ctrl.o_ibus_adr[28] ),
    .A4(_03637_),
    .ZN(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09425_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_adr[30] ),
    .A2(_03561_),
    .B1(_03656_),
    .B2(_03657_),
    .C(_03409_),
    .ZN(_03658_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09426_ (.A1(_03654_),
    .A2(_03658_),
    .ZN(_00072_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09427_ (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[31] ),
    .ZN(_03659_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09428_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[31] ),
    .A2(_03657_),
    .Z(_03660_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09429_ (.A1(_03417_),
    .A2(\mod.u_scanchain_local.module_data_in[68] ),
    .ZN(_03661_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09430_ (.A1(_03659_),
    .A2(_03402_),
    .B1(_03493_),
    .B2(_03660_),
    .C(_03661_),
    .ZN(_00073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09431_ (.I(\mod.u_cpu.cpu.immdec.imm11_7[3] ),
    .Z(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09432_ (.I(_03662_),
    .Z(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09433_ (.I(\mod.u_cpu.cpu.immdec.imm11_7[2] ),
    .Z(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09434_ (.I(\mod.u_cpu.cpu.immdec.imm11_7[4] ),
    .Z(_03665_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _09435_ (.A1(\mod.u_cpu.cpu.immdec.imm11_7[0] ),
    .A2(\mod.u_cpu.cpu.immdec.imm11_7[1] ),
    .A3(_03664_),
    .A4(_03665_),
    .Z(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09436_ (.A1(\mod.u_cpu.cpu.state.init_done ),
    .A2(_01434_),
    .ZN(_03667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09437_ (.A1(_03289_),
    .A2(_03667_),
    .ZN(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09438_ (.I(_03668_),
    .Z(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09439_ (.I(_03331_),
    .Z(_03670_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09440_ (.A1(_03395_),
    .A2(_03331_),
    .ZN(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09441_ (.A1(_03670_),
    .A2(_03403_),
    .B(_03671_),
    .C(_03252_),
    .ZN(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09442_ (.A1(_03663_),
    .A2(_03666_),
    .B(_03669_),
    .C(_03672_),
    .ZN(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09443_ (.I(_03391_),
    .Z(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09444_ (.A1(_03353_),
    .A2(_03673_),
    .B(_03674_),
    .ZN(\mod.u_cpu.cpu.o_wen0 ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09445_ (.A1(_01451_),
    .A2(_03674_),
    .ZN(\mod.u_cpu.cpu.o_wen1 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09446_ (.A1(_03371_),
    .A2(\mod.u_cpu.cpu.ctrl.pc_plus_4_cy_r ),
    .ZN(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09447_ (.A1(_03323_),
    .A2(_03324_),
    .ZN(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09448_ (.A1(_03334_),
    .A2(_03668_),
    .ZN(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09449_ (.A1(_03675_),
    .A2(_03676_),
    .B(_03677_),
    .ZN(_00005_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09450_ (.A1(\mod.u_arbiter.i_wb_cpu_ibus_adr[0] ),
    .A2(\mod.u_cpu.cpu.ctrl.pc_plus_offset_cy_r ),
    .A3(_03265_),
    .ZN(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09451_ (.A1(_03678_),
    .A2(_03294_),
    .B(_03677_),
    .ZN(_00006_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09452_ (.I(\mod.u_cpu.cpu.decode.opcode[1] ),
    .Z(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09453_ (.A1(_03395_),
    .A2(_03679_),
    .ZN(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09454_ (.I(_03255_),
    .Z(_03681_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09455_ (.A1(_03349_),
    .A2(_03681_),
    .ZN(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09456_ (.A1(_03365_),
    .A2(\mod.u_cpu.cpu.bufreg.c_r ),
    .A3(_03680_),
    .A4(_03682_),
    .ZN(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09457_ (.A1(_03356_),
    .A2(_03680_),
    .A3(_03682_),
    .ZN(_03684_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09458_ (.A1(\mod.u_cpu.cpu.bufreg.c_r ),
    .A2(_03684_),
    .ZN(_03685_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09459_ (.I(_03395_),
    .Z(_03686_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09460_ (.A1(_03388_),
    .A2(_03337_),
    .Z(_03687_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09461_ (.A1(_03681_),
    .A2(_03679_),
    .Z(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09462_ (.A1(_03686_),
    .A2(_03687_),
    .A3(_03688_),
    .ZN(_03689_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09463_ (.A1(_03252_),
    .A2(_03276_),
    .A3(_03689_),
    .Z(_03690_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09464_ (.A1(_03685_),
    .A2(_03690_),
    .ZN(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09465_ (.I(_03292_),
    .Z(_03692_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09466_ (.I(_03692_),
    .ZN(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09467_ (.I(_03693_),
    .Z(_03694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09468_ (.A1(_03683_),
    .A2(_03691_),
    .B(_03694_),
    .ZN(_00004_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09469_ (.I0(\mod.u_cpu.rf_ram_if.wdata1_r[0] ),
    .I1(\mod.u_cpu.rf_ram_if.wdata0_r ),
    .S(_01449_),
    .Z(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09470_ (.I(_03695_),
    .Z(_03696_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09471_ (.I(_03696_),
    .Z(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09472_ (.I(_03697_),
    .Z(_03698_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09473_ (.I(_03698_),
    .Z(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09474_ (.A1(_01418_),
    .A2(_01645_),
    .Z(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09475_ (.A1(_01500_),
    .A2(_03700_),
    .ZN(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09476_ (.I(_03701_),
    .Z(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09477_ (.A1(_01439_),
    .A2(_01494_),
    .B(\mod.u_cpu.raddr[1] ),
    .ZN(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09478_ (.A1(_01660_),
    .A2(_03703_),
    .Z(_03704_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09479_ (.A1(\mod.u_cpu.cpu.decode.op21 ),
    .A2(_01426_),
    .B(_01440_),
    .ZN(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09480_ (.A1(_01461_),
    .A2(_03705_),
    .ZN(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09481_ (.A1(\mod.u_cpu.cpu.immdec.imm11_7[0] ),
    .A2(_01441_),
    .B(_03706_),
    .ZN(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09482_ (.A1(_01659_),
    .A2(_03703_),
    .ZN(_03708_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09483_ (.A1(_01531_),
    .A2(_03708_),
    .Z(_03709_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09484_ (.A1(_03707_),
    .A2(_03709_),
    .Z(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09485_ (.A1(_03704_),
    .A2(_03710_),
    .ZN(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09486_ (.A1(_03702_),
    .A2(_03711_),
    .Z(_03712_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09487_ (.I(_03712_),
    .Z(_03713_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09488_ (.I(_03713_),
    .Z(_03714_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09489_ (.A1(_01460_),
    .A2(_03374_),
    .ZN(_03715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09490_ (.A1(_03664_),
    .A2(_03715_),
    .ZN(_03716_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09491_ (.I0(\mod.u_cpu.rf_ram_if.wen1_r ),
    .I1(\mod.u_cpu.rf_ram_if.wen0_r ),
    .S(_01418_),
    .Z(_03717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09492_ (.A1(_03716_),
    .A2(_03717_),
    .ZN(_03718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09493_ (.A1(_01448_),
    .A2(\mod.u_cpu.cpu.immdec.imm11_7[1] ),
    .ZN(_03719_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09494_ (.A1(_01448_),
    .A2(_01454_),
    .B(_03719_),
    .ZN(_03720_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09495_ (.A1(_03374_),
    .A2(_03720_),
    .Z(_03721_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09496_ (.A1(_03718_),
    .A2(_03721_),
    .ZN(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09497_ (.I(_03722_),
    .Z(_03723_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09498_ (.I(_01441_),
    .Z(_03724_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09499_ (.A1(\mod.u_cpu.cpu.immdec.imm11_7[3] ),
    .A2(\mod.u_cpu.cpu.immdec.imm11_7[4] ),
    .A3(_03724_),
    .ZN(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09500_ (.I(_03725_),
    .Z(_03726_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09501_ (.I(_03726_),
    .Z(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09502_ (.A1(_03723_),
    .A2(_03727_),
    .ZN(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09503_ (.A1(_03714_),
    .A2(_03728_),
    .ZN(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09504_ (.I0(\mod.u_cpu.rf_ram.memory[9][0] ),
    .I1(_03699_),
    .S(_03729_),
    .Z(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09505_ (.I(_03730_),
    .Z(_00078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09506_ (.A1(_01462_),
    .A2(\mod.u_cpu.rf_ram_if.wdata1_r[1] ),
    .ZN(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09507_ (.A1(_01462_),
    .A2(_03352_),
    .B(_03731_),
    .ZN(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09508_ (.I(_03732_),
    .Z(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09509_ (.I(_03733_),
    .Z(_03734_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09510_ (.I(_03734_),
    .Z(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09511_ (.I0(\mod.u_cpu.rf_ram.memory[9][1] ),
    .I1(_03735_),
    .S(_03729_),
    .Z(_03736_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09512_ (.I(_03736_),
    .Z(_00079_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09513_ (.I(_03695_),
    .Z(_03737_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09514_ (.I(_03737_),
    .Z(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09515_ (.I(_03738_),
    .Z(_03739_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09516_ (.I(_03739_),
    .Z(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09517_ (.A1(_01461_),
    .A2(_01778_),
    .Z(_03741_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09518_ (.A1(_01418_),
    .A2(_01498_),
    .A3(_01518_),
    .Z(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09519_ (.A1(_03703_),
    .A2(_03742_),
    .Z(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09520_ (.A1(_03741_),
    .A2(_03743_),
    .ZN(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09521_ (.I(_03744_),
    .Z(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09522_ (.A1(_01850_),
    .A2(_03703_),
    .Z(_03746_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09523_ (.A1(_03271_),
    .A2(_03715_),
    .B1(_03705_),
    .B2(_01461_),
    .ZN(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09524_ (.I(_03709_),
    .Z(_03748_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09525_ (.A1(_03746_),
    .A2(_03747_),
    .A3(_03748_),
    .ZN(_03749_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09526_ (.A1(_03745_),
    .A2(_03749_),
    .ZN(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09527_ (.I(_03750_),
    .Z(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09528_ (.I(_03751_),
    .Z(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09529_ (.I(_03715_),
    .Z(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09530_ (.A1(_03716_),
    .A2(_03717_),
    .Z(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09531_ (.A1(_03754_),
    .A2(_03721_),
    .ZN(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09532_ (.A1(_03753_),
    .A2(_03755_),
    .ZN(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09533_ (.I(_03756_),
    .Z(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09534_ (.I(_03757_),
    .Z(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09535_ (.A1(_03752_),
    .A2(_03758_),
    .ZN(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09536_ (.I0(_03740_),
    .I1(\mod.u_cpu.rf_ram.memory[574][0] ),
    .S(_03759_),
    .Z(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09537_ (.I(_03760_),
    .Z(_00080_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09538_ (.I(_03732_),
    .Z(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09539_ (.I(_03761_),
    .Z(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09540_ (.I(_03762_),
    .Z(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09541_ (.I(_03763_),
    .Z(_03764_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09542_ (.I0(_03764_),
    .I1(\mod.u_cpu.rf_ram.memory[574][1] ),
    .S(_03759_),
    .Z(_03765_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09543_ (.I(_03765_),
    .Z(_00081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09544_ (.I(_03756_),
    .Z(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09545_ (.I(_03766_),
    .Z(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09546_ (.I(_03701_),
    .Z(_03768_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09547_ (.A1(_03768_),
    .A2(_03749_),
    .ZN(_03769_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09548_ (.I(_03769_),
    .Z(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09549_ (.I(_03770_),
    .Z(_03771_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09550_ (.A1(_03767_),
    .A2(_03771_),
    .ZN(_03772_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09551_ (.I(_03695_),
    .Z(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09552_ (.I(_03773_),
    .Z(_03774_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09553_ (.I(_03774_),
    .Z(_03775_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09554_ (.A1(_03775_),
    .A2(_03772_),
    .ZN(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09555_ (.A1(_02497_),
    .A2(_03772_),
    .B(_03776_),
    .ZN(_00082_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09556_ (.I0(_03764_),
    .I1(\mod.u_cpu.rf_ram.memory[573][1] ),
    .S(_03772_),
    .Z(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09557_ (.I(_03777_),
    .Z(_00083_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09558_ (.A1(_03700_),
    .A2(_03743_),
    .Z(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09559_ (.I(_03778_),
    .Z(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09560_ (.A1(_03749_),
    .A2(_03779_),
    .ZN(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09561_ (.I(_03780_),
    .Z(_03781_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09562_ (.I(_03781_),
    .Z(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09563_ (.A1(_03758_),
    .A2(_03782_),
    .ZN(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09564_ (.I0(_03740_),
    .I1(\mod.u_cpu.rf_ram.memory[572][0] ),
    .S(_03783_),
    .Z(_03784_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09565_ (.I(_03784_),
    .Z(_00084_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09566_ (.I0(_03764_),
    .I1(\mod.u_cpu.rf_ram.memory[572][1] ),
    .S(_03783_),
    .Z(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09567_ (.I(_03785_),
    .Z(_00085_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09568_ (.A1(_03704_),
    .A2(_03747_),
    .A3(_03748_),
    .ZN(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09569_ (.A1(_03700_),
    .A2(_03743_),
    .ZN(_03787_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09570_ (.I(_03787_),
    .Z(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09571_ (.A1(_03786_),
    .A2(_03788_),
    .ZN(_03789_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09572_ (.I(_03789_),
    .Z(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09573_ (.I(_03790_),
    .Z(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09574_ (.A1(_03758_),
    .A2(_03791_),
    .ZN(_03792_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09575_ (.I0(_03740_),
    .I1(\mod.u_cpu.rf_ram.memory[571][0] ),
    .S(_03792_),
    .Z(_03793_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09576_ (.I(_03793_),
    .Z(_00086_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09577_ (.I0(_03764_),
    .I1(\mod.u_cpu.rf_ram.memory[571][1] ),
    .S(_03792_),
    .Z(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09578_ (.I(_03794_),
    .Z(_00087_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09579_ (.A1(_03745_),
    .A2(_03786_),
    .ZN(_03795_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09580_ (.I(_03795_),
    .Z(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09581_ (.I(_03796_),
    .Z(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09582_ (.A1(_03758_),
    .A2(_03797_),
    .ZN(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09583_ (.I0(_03740_),
    .I1(\mod.u_cpu.rf_ram.memory[570][0] ),
    .S(_03798_),
    .Z(_03799_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09584_ (.I(_03799_),
    .Z(_00088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09585_ (.I(_03763_),
    .Z(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09586_ (.I0(_03800_),
    .I1(\mod.u_cpu.rf_ram.memory[570][1] ),
    .S(_03798_),
    .Z(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09587_ (.I(_03801_),
    .Z(_00089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09588_ (.I(_03739_),
    .Z(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09589_ (.A1(_03779_),
    .A2(_03786_),
    .ZN(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09590_ (.I(_03803_),
    .Z(_03804_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09591_ (.I(_03804_),
    .Z(_03805_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09592_ (.A1(_03374_),
    .A2(_03720_),
    .ZN(_03806_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09593_ (.A1(_03718_),
    .A2(_03806_),
    .ZN(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09594_ (.A1(_03725_),
    .A2(_03807_),
    .Z(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09595_ (.I(_03808_),
    .Z(_03809_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09596_ (.I(_03809_),
    .Z(_03810_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09597_ (.A1(_03805_),
    .A2(_03810_),
    .ZN(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09598_ (.I0(_03802_),
    .I1(\mod.u_cpu.rf_ram.memory[56][0] ),
    .S(_03811_),
    .Z(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09599_ (.I(_03812_),
    .Z(_00090_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09600_ (.I0(_03800_),
    .I1(\mod.u_cpu.rf_ram.memory[56][1] ),
    .S(_03811_),
    .Z(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09601_ (.I(_03813_),
    .Z(_00091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09602_ (.I(_03757_),
    .Z(_03814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09603_ (.A1(_03814_),
    .A2(_03805_),
    .ZN(_03815_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09604_ (.I0(_03802_),
    .I1(\mod.u_cpu.rf_ram.memory[568][0] ),
    .S(_03815_),
    .Z(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09605_ (.I(_03816_),
    .Z(_00092_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09606_ (.I0(_03800_),
    .I1(\mod.u_cpu.rf_ram.memory[568][1] ),
    .S(_03815_),
    .Z(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09607_ (.I(_03817_),
    .Z(_00093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09608_ (.I(_03787_),
    .Z(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09609_ (.A1(_03707_),
    .A2(_03748_),
    .ZN(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09610_ (.A1(_03746_),
    .A2(_03819_),
    .ZN(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09611_ (.A1(_03818_),
    .A2(_03820_),
    .ZN(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09612_ (.I(_03821_),
    .Z(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09613_ (.I(_03822_),
    .Z(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09614_ (.A1(_03767_),
    .A2(_03823_),
    .ZN(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09615_ (.A1(_03775_),
    .A2(_03824_),
    .ZN(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09616_ (.A1(_02513_),
    .A2(_03824_),
    .B(_03825_),
    .ZN(_00094_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09617_ (.I0(_03800_),
    .I1(\mod.u_cpu.rf_ram.memory[567][1] ),
    .S(_03824_),
    .Z(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09618_ (.I(_03826_),
    .Z(_00095_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09619_ (.A1(_03745_),
    .A2(_03820_),
    .ZN(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09620_ (.I(_03827_),
    .Z(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09621_ (.I(_03828_),
    .Z(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09622_ (.A1(_03814_),
    .A2(_03829_),
    .ZN(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09623_ (.I0(_03802_),
    .I1(\mod.u_cpu.rf_ram.memory[566][0] ),
    .S(_03830_),
    .Z(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09624_ (.I(_03831_),
    .Z(_00096_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09625_ (.I(_03763_),
    .Z(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09626_ (.I0(_03832_),
    .I1(\mod.u_cpu.rf_ram.memory[566][1] ),
    .S(_03830_),
    .Z(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09627_ (.I(_03833_),
    .Z(_00097_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09628_ (.I(_03766_),
    .Z(_03834_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09629_ (.A1(_03702_),
    .A2(_03820_),
    .ZN(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09630_ (.I(_03835_),
    .Z(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09631_ (.I(_03836_),
    .Z(_03837_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09632_ (.A1(_03834_),
    .A2(_03837_),
    .ZN(_03838_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09633_ (.A1(_03775_),
    .A2(_03838_),
    .ZN(_03839_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09634_ (.A1(_02510_),
    .A2(_03838_),
    .B(_03839_),
    .ZN(_00098_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09635_ (.I0(_03832_),
    .I1(\mod.u_cpu.rf_ram.memory[565][1] ),
    .S(_03838_),
    .Z(_03840_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09636_ (.I(_03840_),
    .Z(_00099_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09637_ (.A1(_03779_),
    .A2(_03820_),
    .ZN(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09638_ (.I(_03841_),
    .Z(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09639_ (.I(_03842_),
    .Z(_03843_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09640_ (.A1(_03814_),
    .A2(_03843_),
    .ZN(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09641_ (.I0(_03802_),
    .I1(\mod.u_cpu.rf_ram.memory[564][0] ),
    .S(_03844_),
    .Z(_03845_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09642_ (.I(_03845_),
    .Z(_00100_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09643_ (.I0(_03832_),
    .I1(\mod.u_cpu.rf_ram.memory[564][1] ),
    .S(_03844_),
    .Z(_03846_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09644_ (.I(_03846_),
    .Z(_00101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09645_ (.I(_03739_),
    .Z(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09646_ (.A1(_03704_),
    .A2(_03819_),
    .ZN(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09647_ (.A1(_03788_),
    .A2(_03848_),
    .ZN(_03849_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09648_ (.I(_03849_),
    .Z(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09649_ (.I(_03850_),
    .Z(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09650_ (.A1(_03814_),
    .A2(_03851_),
    .ZN(_03852_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09651_ (.I0(_03847_),
    .I1(\mod.u_cpu.rf_ram.memory[563][0] ),
    .S(_03852_),
    .Z(_03853_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09652_ (.I(_03853_),
    .Z(_00102_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09653_ (.I0(_03832_),
    .I1(\mod.u_cpu.rf_ram.memory[563][1] ),
    .S(_03852_),
    .Z(_03854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09654_ (.I(_03854_),
    .Z(_00103_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09655_ (.I(_03757_),
    .Z(_03855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09656_ (.I(_03744_),
    .Z(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09657_ (.A1(_03856_),
    .A2(_03848_),
    .ZN(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09658_ (.I(_03857_),
    .Z(_03858_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09659_ (.I(_03858_),
    .Z(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09660_ (.A1(_03855_),
    .A2(_03859_),
    .ZN(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09661_ (.I0(_03847_),
    .I1(\mod.u_cpu.rf_ram.memory[562][0] ),
    .S(_03860_),
    .Z(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09662_ (.I(_03861_),
    .Z(_00104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09663_ (.I(_03763_),
    .Z(_03862_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09664_ (.I0(_03862_),
    .I1(\mod.u_cpu.rf_ram.memory[562][1] ),
    .S(_03860_),
    .Z(_03863_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09665_ (.I(_03863_),
    .Z(_00105_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09666_ (.A1(_03768_),
    .A2(_03848_),
    .ZN(_03864_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09667_ (.I(_03864_),
    .Z(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09668_ (.I(_03865_),
    .Z(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09669_ (.A1(_03855_),
    .A2(_03866_),
    .ZN(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09670_ (.I0(_03847_),
    .I1(\mod.u_cpu.rf_ram.memory[561][0] ),
    .S(_03867_),
    .Z(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09671_ (.I(_03868_),
    .Z(_00106_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09672_ (.I0(_03862_),
    .I1(\mod.u_cpu.rf_ram.memory[561][1] ),
    .S(_03867_),
    .Z(_03869_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09673_ (.I(_03869_),
    .Z(_00107_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09674_ (.I(_03778_),
    .Z(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09675_ (.A1(_03870_),
    .A2(_03848_),
    .ZN(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09676_ (.I(_03871_),
    .Z(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09677_ (.I(_03872_),
    .Z(_03873_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09678_ (.A1(_03855_),
    .A2(_03873_),
    .ZN(_03874_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09679_ (.I0(_03847_),
    .I1(\mod.u_cpu.rf_ram.memory[560][0] ),
    .S(_03874_),
    .Z(_03875_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09680_ (.I(_03875_),
    .Z(_00108_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09681_ (.I0(_03862_),
    .I1(\mod.u_cpu.rf_ram.memory[560][1] ),
    .S(_03874_),
    .Z(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09682_ (.I(_03876_),
    .Z(_00109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09683_ (.I(_03739_),
    .Z(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09684_ (.I(_03809_),
    .Z(_03878_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09685_ (.I(_03822_),
    .Z(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09686_ (.A1(_03878_),
    .A2(_03879_),
    .ZN(_03880_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09687_ (.I0(_03877_),
    .I1(\mod.u_cpu.rf_ram.memory[55][0] ),
    .S(_03880_),
    .Z(_03881_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09688_ (.I(_03881_),
    .Z(_00110_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09689_ (.I0(_03862_),
    .I1(\mod.u_cpu.rf_ram.memory[55][1] ),
    .S(_03880_),
    .Z(_03882_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09690_ (.I(_03882_),
    .Z(_00111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09691_ (.A1(_03746_),
    .A2(_03710_),
    .ZN(_03883_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09692_ (.A1(_03856_),
    .A2(_03883_),
    .ZN(_03884_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09693_ (.I(_03884_),
    .Z(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09694_ (.I(_03885_),
    .Z(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09695_ (.A1(_03855_),
    .A2(_03886_),
    .ZN(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09696_ (.I0(_03877_),
    .I1(\mod.u_cpu.rf_ram.memory[558][0] ),
    .S(_03887_),
    .Z(_03888_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09697_ (.I(_03888_),
    .Z(_00112_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09698_ (.I(_03762_),
    .Z(_03889_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09699_ (.I(_03889_),
    .Z(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09700_ (.I0(_03890_),
    .I1(\mod.u_cpu.rf_ram.memory[558][1] ),
    .S(_03887_),
    .Z(_03891_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09701_ (.I(_03891_),
    .Z(_00113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09702_ (.I(_03807_),
    .Z(_03892_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09703_ (.A1(_03724_),
    .A2(_03892_),
    .ZN(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09704_ (.A1(_03702_),
    .A2(_03883_),
    .Z(_03894_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09705_ (.I(_03894_),
    .Z(_03895_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09706_ (.I(_03895_),
    .Z(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09707_ (.A1(_03893_),
    .A2(_03896_),
    .ZN(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09708_ (.I(_03697_),
    .Z(_03898_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09709_ (.I(_03898_),
    .Z(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09710_ (.A1(_03899_),
    .A2(_03897_),
    .ZN(_03900_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09711_ (.A1(_02480_),
    .A2(_03897_),
    .B(_03900_),
    .ZN(_00114_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09712_ (.I0(\mod.u_cpu.rf_ram.memory[557][1] ),
    .I1(_03735_),
    .S(_03897_),
    .Z(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09713_ (.I(_03901_),
    .Z(_00115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09714_ (.I(_03766_),
    .Z(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09715_ (.A1(_03870_),
    .A2(_03883_),
    .ZN(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09716_ (.I(_03903_),
    .Z(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09717_ (.I(_03904_),
    .Z(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09718_ (.A1(_03902_),
    .A2(_03905_),
    .ZN(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09719_ (.I0(_03877_),
    .I1(\mod.u_cpu.rf_ram.memory[556][0] ),
    .S(_03906_),
    .Z(_03907_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09720_ (.I(_03907_),
    .Z(_00116_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09721_ (.I0(_03890_),
    .I1(\mod.u_cpu.rf_ram.memory[556][1] ),
    .S(_03906_),
    .Z(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09722_ (.I(_03908_),
    .Z(_00117_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09723_ (.A1(_03711_),
    .A2(_03788_),
    .ZN(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09724_ (.I(_03909_),
    .Z(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09725_ (.I(_03910_),
    .Z(_03911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09726_ (.A1(_03902_),
    .A2(_03911_),
    .ZN(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09727_ (.I0(_03877_),
    .I1(\mod.u_cpu.rf_ram.memory[555][0] ),
    .S(_03912_),
    .Z(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09728_ (.I(_03913_),
    .Z(_00118_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09729_ (.I0(_03890_),
    .I1(\mod.u_cpu.rf_ram.memory[555][1] ),
    .S(_03912_),
    .Z(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09730_ (.I(_03914_),
    .Z(_00119_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09731_ (.I(_03738_),
    .Z(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09732_ (.I(_03915_),
    .Z(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09733_ (.A1(_03711_),
    .A2(_03745_),
    .ZN(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09734_ (.I(_03917_),
    .Z(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09735_ (.I(_03918_),
    .Z(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09736_ (.A1(_03902_),
    .A2(_03919_),
    .ZN(_03920_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09737_ (.I0(_03916_),
    .I1(\mod.u_cpu.rf_ram.memory[554][0] ),
    .S(_03920_),
    .Z(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09738_ (.I(_03921_),
    .Z(_00120_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09739_ (.I0(_03890_),
    .I1(\mod.u_cpu.rf_ram.memory[554][1] ),
    .S(_03920_),
    .Z(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09740_ (.I(_03922_),
    .Z(_00121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09741_ (.I(_03696_),
    .Z(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09742_ (.I(_03923_),
    .Z(_03924_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09743_ (.I(_03924_),
    .Z(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09744_ (.A1(_03714_),
    .A2(_03893_),
    .ZN(_03926_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09745_ (.I0(\mod.u_cpu.rf_ram.memory[553][0] ),
    .I1(_03925_),
    .S(_03926_),
    .Z(_03927_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09746_ (.I(_03927_),
    .Z(_00122_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09747_ (.I(_03733_),
    .Z(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09748_ (.I(_03928_),
    .Z(_03929_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09749_ (.I0(\mod.u_cpu.rf_ram.memory[553][1] ),
    .I1(_03929_),
    .S(_03926_),
    .Z(_03930_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09750_ (.I(_03930_),
    .Z(_00123_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09751_ (.A1(_03711_),
    .A2(_03779_),
    .ZN(_03931_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09752_ (.I(_03931_),
    .Z(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09753_ (.I(_03932_),
    .Z(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09754_ (.A1(_03902_),
    .A2(_03933_),
    .ZN(_03934_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09755_ (.I0(_03916_),
    .I1(\mod.u_cpu.rf_ram.memory[552][0] ),
    .S(_03934_),
    .Z(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09756_ (.I(_03935_),
    .Z(_00124_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09757_ (.I(_03889_),
    .Z(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09758_ (.I0(_03936_),
    .I1(\mod.u_cpu.rf_ram.memory[552][1] ),
    .S(_03934_),
    .Z(_03937_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09759_ (.I(_03937_),
    .Z(_00125_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09760_ (.A1(_03747_),
    .A2(_03748_),
    .ZN(_03938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09761_ (.A1(_03746_),
    .A2(_03938_),
    .ZN(_03939_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09762_ (.A1(_03818_),
    .A2(_03939_),
    .ZN(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09763_ (.I(_03940_),
    .Z(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09764_ (.I(_03941_),
    .Z(_03942_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09765_ (.A1(_03834_),
    .A2(_03942_),
    .ZN(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09766_ (.I(_03697_),
    .Z(_03944_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09767_ (.I(_03944_),
    .Z(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09768_ (.A1(_03945_),
    .A2(_03943_),
    .ZN(_03946_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09769_ (.A1(_02463_),
    .A2(_03943_),
    .B(_03946_),
    .ZN(_00126_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09770_ (.I0(_03936_),
    .I1(\mod.u_cpu.rf_ram.memory[551][1] ),
    .S(_03943_),
    .Z(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09771_ (.I(_03947_),
    .Z(_00127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09772_ (.I(_03766_),
    .Z(_03948_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09773_ (.A1(_03856_),
    .A2(_03939_),
    .ZN(_03949_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09774_ (.I(_03949_),
    .Z(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09775_ (.I(_03950_),
    .Z(_03951_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09776_ (.A1(_03948_),
    .A2(_03951_),
    .ZN(_03952_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09777_ (.I0(_03916_),
    .I1(\mod.u_cpu.rf_ram.memory[550][0] ),
    .S(_03952_),
    .Z(_03953_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09778_ (.I(_03953_),
    .Z(_00128_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09779_ (.I0(_03936_),
    .I1(\mod.u_cpu.rf_ram.memory[550][1] ),
    .S(_03952_),
    .Z(_03954_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09780_ (.I(_03954_),
    .Z(_00129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09781_ (.A1(_03878_),
    .A2(_03829_),
    .ZN(_03955_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09782_ (.I0(_03916_),
    .I1(\mod.u_cpu.rf_ram.memory[54][0] ),
    .S(_03955_),
    .Z(_03956_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09783_ (.I(_03956_),
    .Z(_00130_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09784_ (.I0(_03936_),
    .I1(\mod.u_cpu.rf_ram.memory[54][1] ),
    .S(_03955_),
    .Z(_03957_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09785_ (.I(_03957_),
    .Z(_00131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09786_ (.I(_03915_),
    .Z(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09787_ (.A1(_03870_),
    .A2(_03939_),
    .ZN(_03959_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09788_ (.I(_03959_),
    .Z(_03960_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09789_ (.I(_03960_),
    .Z(_03961_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09790_ (.A1(_03948_),
    .A2(_03961_),
    .ZN(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09791_ (.I0(_03958_),
    .I1(\mod.u_cpu.rf_ram.memory[548][0] ),
    .S(_03962_),
    .Z(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09792_ (.I(_03963_),
    .Z(_00132_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09793_ (.I(_03889_),
    .Z(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09794_ (.I0(_03964_),
    .I1(\mod.u_cpu.rf_ram.memory[548][1] ),
    .S(_03962_),
    .Z(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09795_ (.I(_03965_),
    .Z(_00133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09796_ (.A1(_03704_),
    .A2(_03938_),
    .ZN(_03966_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09797_ (.A1(_03788_),
    .A2(_03966_),
    .ZN(_03967_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09798_ (.I(_03967_),
    .Z(_03968_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09799_ (.I(_03968_),
    .Z(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09800_ (.A1(_03948_),
    .A2(_03969_),
    .ZN(_03970_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09801_ (.I0(_03958_),
    .I1(\mod.u_cpu.rf_ram.memory[547][0] ),
    .S(_03970_),
    .Z(_03971_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09802_ (.I(_03971_),
    .Z(_00134_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09803_ (.I0(_03964_),
    .I1(\mod.u_cpu.rf_ram.memory[547][1] ),
    .S(_03970_),
    .Z(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09804_ (.I(_03972_),
    .Z(_00135_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09805_ (.A1(_03856_),
    .A2(_03966_),
    .ZN(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09806_ (.I(_03973_),
    .Z(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09807_ (.I(_03974_),
    .Z(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09808_ (.A1(_03948_),
    .A2(_03975_),
    .ZN(_03976_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09809_ (.I0(_03958_),
    .I1(\mod.u_cpu.rf_ram.memory[546][0] ),
    .S(_03976_),
    .Z(_03977_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09810_ (.I(_03977_),
    .Z(_00136_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09811_ (.I0(_03964_),
    .I1(\mod.u_cpu.rf_ram.memory[546][1] ),
    .S(_03976_),
    .Z(_03978_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09812_ (.I(_03978_),
    .Z(_00137_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09813_ (.A1(_03768_),
    .A2(_03966_),
    .ZN(_03979_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09814_ (.I(_03979_),
    .Z(_03980_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09815_ (.A1(_03757_),
    .A2(_03980_),
    .Z(_03981_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09816_ (.I0(\mod.u_cpu.rf_ram.memory[545][0] ),
    .I1(_03925_),
    .S(_03981_),
    .Z(_03982_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09817_ (.I(_03982_),
    .Z(_00138_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09818_ (.I0(\mod.u_cpu.rf_ram.memory[545][1] ),
    .I1(_03929_),
    .S(_03981_),
    .Z(_03983_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09819_ (.I(_03983_),
    .Z(_00139_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09820_ (.A1(_03870_),
    .A2(_03966_),
    .ZN(_03984_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09821_ (.I(_03984_),
    .Z(_03985_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09822_ (.I(_03985_),
    .Z(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09823_ (.A1(_03767_),
    .A2(_03986_),
    .ZN(_03987_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09824_ (.I0(_03958_),
    .I1(\mod.u_cpu.rf_ram.memory[544][0] ),
    .S(_03987_),
    .Z(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09825_ (.I(_03988_),
    .Z(_00140_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09826_ (.I0(_03964_),
    .I1(\mod.u_cpu.rf_ram.memory[544][1] ),
    .S(_03987_),
    .Z(_03989_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09827_ (.I(_03989_),
    .Z(_00141_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09828_ (.A1(_03749_),
    .A2(_03818_),
    .ZN(_03990_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09829_ (.I(_03990_),
    .Z(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09830_ (.I(_03806_),
    .Z(_03992_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09831_ (.A1(_03754_),
    .A2(_03992_),
    .ZN(_03993_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09832_ (.A1(_01478_),
    .A2(_03993_),
    .ZN(_03994_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09833_ (.I(_03994_),
    .Z(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09834_ (.I(_03995_),
    .Z(_03996_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09835_ (.A1(_03991_),
    .A2(_03996_),
    .ZN(_03997_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09836_ (.A1(_03945_),
    .A2(_03997_),
    .ZN(_03998_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09837_ (.A1(_02576_),
    .A2(_03997_),
    .B(_03998_),
    .ZN(_00142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09838_ (.I(_03889_),
    .Z(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09839_ (.I0(_03999_),
    .I1(\mod.u_cpu.rf_ram.memory[543][1] ),
    .S(_03997_),
    .Z(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09840_ (.I(_04000_),
    .Z(_00143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09841_ (.I(_03915_),
    .Z(_04001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09842_ (.I(_03994_),
    .Z(_04002_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09843_ (.I(_04002_),
    .Z(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09844_ (.A1(_03752_),
    .A2(_04003_),
    .ZN(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09845_ (.I0(_04001_),
    .I1(\mod.u_cpu.rf_ram.memory[542][0] ),
    .S(_04004_),
    .Z(_04005_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09846_ (.I(_04005_),
    .Z(_00144_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09847_ (.I0(_03999_),
    .I1(\mod.u_cpu.rf_ram.memory[542][1] ),
    .S(_04004_),
    .Z(_04006_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09848_ (.I(_04006_),
    .Z(_00145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09849_ (.A1(_03771_),
    .A2(_03996_),
    .ZN(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09850_ (.A1(_03945_),
    .A2(_04007_),
    .ZN(_04008_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09851_ (.A1(_02573_),
    .A2(_04007_),
    .B(_04008_),
    .ZN(_00146_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09852_ (.I0(_03999_),
    .I1(\mod.u_cpu.rf_ram.memory[541][1] ),
    .S(_04007_),
    .Z(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09853_ (.I(_04009_),
    .Z(_00147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09854_ (.A1(_03782_),
    .A2(_04003_),
    .ZN(_04010_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09855_ (.I0(_04001_),
    .I1(\mod.u_cpu.rf_ram.memory[540][0] ),
    .S(_04010_),
    .Z(_04011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09856_ (.I(_04011_),
    .Z(_00148_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09857_ (.I0(_03999_),
    .I1(\mod.u_cpu.rf_ram.memory[540][1] ),
    .S(_04010_),
    .Z(_04012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09858_ (.I(_04012_),
    .Z(_00149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09859_ (.I(_03809_),
    .Z(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09860_ (.I(_03836_),
    .Z(_04014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09861_ (.A1(_04013_),
    .A2(_04014_),
    .ZN(_04015_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09862_ (.I0(_04001_),
    .I1(\mod.u_cpu.rf_ram.memory[53][0] ),
    .S(_04015_),
    .Z(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09863_ (.I(_04016_),
    .Z(_00150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09864_ (.I(_03762_),
    .Z(_04017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09865_ (.I(_04017_),
    .Z(_04018_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09866_ (.I0(_04018_),
    .I1(\mod.u_cpu.rf_ram.memory[53][1] ),
    .S(_04015_),
    .Z(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09867_ (.I(_04019_),
    .Z(_00151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09868_ (.A1(_03797_),
    .A2(_04003_),
    .ZN(_04020_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09869_ (.I0(_04001_),
    .I1(\mod.u_cpu.rf_ram.memory[538][0] ),
    .S(_04020_),
    .Z(_04021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09870_ (.I(_04021_),
    .Z(_00152_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09871_ (.I0(_04018_),
    .I1(\mod.u_cpu.rf_ram.memory[538][1] ),
    .S(_04020_),
    .Z(_04022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09872_ (.I(_04022_),
    .Z(_00153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09873_ (.I(_03915_),
    .Z(_04023_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09874_ (.A1(_03768_),
    .A2(_03786_),
    .ZN(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09875_ (.I(_04024_),
    .Z(_04025_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09876_ (.I(_04025_),
    .Z(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09877_ (.A1(_03996_),
    .A2(_04026_),
    .ZN(_04027_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09878_ (.I0(_04023_),
    .I1(\mod.u_cpu.rf_ram.memory[537][0] ),
    .S(_04027_),
    .Z(_04028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09879_ (.I(_04028_),
    .Z(_00154_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09880_ (.I0(_04018_),
    .I1(\mod.u_cpu.rf_ram.memory[537][1] ),
    .S(_04027_),
    .Z(_04029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09881_ (.I(_04029_),
    .Z(_00155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09882_ (.A1(_03805_),
    .A2(_04003_),
    .ZN(_04030_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09883_ (.I0(_04023_),
    .I1(\mod.u_cpu.rf_ram.memory[536][0] ),
    .S(_04030_),
    .Z(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09884_ (.I(_04031_),
    .Z(_00156_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09885_ (.I0(_04018_),
    .I1(\mod.u_cpu.rf_ram.memory[536][1] ),
    .S(_04030_),
    .Z(_04032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09886_ (.I(_04032_),
    .Z(_00157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09887_ (.I(_03995_),
    .Z(_04033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09888_ (.A1(_03823_),
    .A2(_04033_),
    .ZN(_04034_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09889_ (.A1(_03945_),
    .A2(_04034_),
    .ZN(_04035_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09890_ (.A1(_02567_),
    .A2(_04034_),
    .B(_04035_),
    .ZN(_00158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09891_ (.I(_04017_),
    .Z(_04036_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09892_ (.I0(_04036_),
    .I1(\mod.u_cpu.rf_ram.memory[535][1] ),
    .S(_04034_),
    .Z(_04037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09893_ (.I(_04037_),
    .Z(_00159_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09894_ (.I(_04002_),
    .Z(_04038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09895_ (.A1(_03829_),
    .A2(_04038_),
    .ZN(_04039_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09896_ (.I0(_04023_),
    .I1(\mod.u_cpu.rf_ram.memory[534][0] ),
    .S(_04039_),
    .Z(_04040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09897_ (.I(_04040_),
    .Z(_00160_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09898_ (.I0(_04036_),
    .I1(\mod.u_cpu.rf_ram.memory[534][1] ),
    .S(_04039_),
    .Z(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09899_ (.I(_04041_),
    .Z(_00161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09900_ (.A1(_03837_),
    .A2(_04033_),
    .ZN(_04042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09901_ (.I(_03697_),
    .Z(_04043_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09902_ (.I(_04043_),
    .Z(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09903_ (.A1(_04044_),
    .A2(_04042_),
    .ZN(_04045_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09904_ (.A1(_02563_),
    .A2(_04042_),
    .B(_04045_),
    .ZN(_00162_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09905_ (.I0(_04036_),
    .I1(\mod.u_cpu.rf_ram.memory[533][1] ),
    .S(_04042_),
    .Z(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09906_ (.I(_04046_),
    .Z(_00163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09907_ (.A1(_03843_),
    .A2(_04038_),
    .ZN(_04047_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09908_ (.I0(_04023_),
    .I1(\mod.u_cpu.rf_ram.memory[532][0] ),
    .S(_04047_),
    .Z(_04048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09909_ (.I(_04048_),
    .Z(_00164_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09910_ (.I0(_04036_),
    .I1(\mod.u_cpu.rf_ram.memory[532][1] ),
    .S(_04047_),
    .Z(_04049_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09911_ (.I(_04049_),
    .Z(_00165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09912_ (.I(_03738_),
    .Z(_04050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09913_ (.I(_04050_),
    .Z(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09914_ (.A1(_03851_),
    .A2(_04038_),
    .ZN(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09915_ (.I0(_04051_),
    .I1(\mod.u_cpu.rf_ram.memory[531][0] ),
    .S(_04052_),
    .Z(_04053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09916_ (.I(_04053_),
    .Z(_00166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09917_ (.I(_04017_),
    .Z(_04054_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09918_ (.I0(_04054_),
    .I1(\mod.u_cpu.rf_ram.memory[531][1] ),
    .S(_04052_),
    .Z(_04055_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09919_ (.I(_04055_),
    .Z(_00167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09920_ (.A1(_03859_),
    .A2(_04038_),
    .ZN(_04056_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09921_ (.I0(_04051_),
    .I1(\mod.u_cpu.rf_ram.memory[530][0] ),
    .S(_04056_),
    .Z(_04057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09922_ (.I(_04057_),
    .Z(_00168_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09923_ (.I0(_04054_),
    .I1(\mod.u_cpu.rf_ram.memory[530][1] ),
    .S(_04056_),
    .Z(_04058_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09924_ (.I(_04058_),
    .Z(_00169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09925_ (.A1(_04013_),
    .A2(_03843_),
    .ZN(_04059_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09926_ (.I0(_04051_),
    .I1(\mod.u_cpu.rf_ram.memory[52][0] ),
    .S(_04059_),
    .Z(_04060_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09927_ (.I(_04060_),
    .Z(_00170_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09928_ (.I0(_04054_),
    .I1(\mod.u_cpu.rf_ram.memory[52][1] ),
    .S(_04059_),
    .Z(_04061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09929_ (.I(_04061_),
    .Z(_00171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09930_ (.I(_04002_),
    .Z(_04062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09931_ (.A1(_03873_),
    .A2(_04062_),
    .ZN(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09932_ (.I0(_04051_),
    .I1(\mod.u_cpu.rf_ram.memory[528][0] ),
    .S(_04063_),
    .Z(_04064_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09933_ (.I(_04064_),
    .Z(_00172_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09934_ (.I0(_04054_),
    .I1(\mod.u_cpu.rf_ram.memory[528][1] ),
    .S(_04063_),
    .Z(_04065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09935_ (.I(_04065_),
    .Z(_00173_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09936_ (.A1(_03818_),
    .A2(_03883_),
    .ZN(_04066_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09937_ (.I(_04066_),
    .Z(_04067_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09938_ (.I(_04067_),
    .Z(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09939_ (.A1(_04033_),
    .A2(_04068_),
    .ZN(_04069_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09940_ (.A1(_04044_),
    .A2(_04069_),
    .ZN(_04070_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09941_ (.A1(_02552_),
    .A2(_04069_),
    .B(_04070_),
    .ZN(_00174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09942_ (.I(_04017_),
    .Z(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09943_ (.I0(_04071_),
    .I1(\mod.u_cpu.rf_ram.memory[527][1] ),
    .S(_04069_),
    .Z(_04072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09944_ (.I(_04072_),
    .Z(_00175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09945_ (.I(_04050_),
    .Z(_04073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09946_ (.A1(_03886_),
    .A2(_04062_),
    .ZN(_04074_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09947_ (.I0(_04073_),
    .I1(\mod.u_cpu.rf_ram.memory[526][0] ),
    .S(_04074_),
    .Z(_04075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09948_ (.I(_04075_),
    .Z(_00176_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09949_ (.I0(_04071_),
    .I1(\mod.u_cpu.rf_ram.memory[526][1] ),
    .S(_04074_),
    .Z(_04076_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09950_ (.I(_04076_),
    .Z(_00177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09951_ (.A1(_01463_),
    .A2(_03722_),
    .ZN(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09952_ (.A1(_03896_),
    .A2(_04077_),
    .ZN(_04078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09953_ (.A1(_03899_),
    .A2(_04078_),
    .ZN(_04079_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09954_ (.A1(_02547_),
    .A2(_04078_),
    .B(_04079_),
    .ZN(_00178_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09955_ (.I0(\mod.u_cpu.rf_ram.memory[525][1] ),
    .I1(_03929_),
    .S(_04078_),
    .Z(_04080_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09956_ (.I(_04080_),
    .Z(_00179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09957_ (.A1(_03905_),
    .A2(_04062_),
    .ZN(_04081_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09958_ (.I0(_04073_),
    .I1(\mod.u_cpu.rf_ram.memory[524][0] ),
    .S(_04081_),
    .Z(_04082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09959_ (.I(_04082_),
    .Z(_00180_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09960_ (.I0(_04071_),
    .I1(\mod.u_cpu.rf_ram.memory[524][1] ),
    .S(_04081_),
    .Z(_04083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09961_ (.I(_04083_),
    .Z(_00181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09962_ (.A1(_03911_),
    .A2(_04062_),
    .ZN(_04084_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09963_ (.I0(_04073_),
    .I1(\mod.u_cpu.rf_ram.memory[523][0] ),
    .S(_04084_),
    .Z(_04085_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09964_ (.I(_04085_),
    .Z(_00182_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09965_ (.I0(_04071_),
    .I1(\mod.u_cpu.rf_ram.memory[523][1] ),
    .S(_04084_),
    .Z(_04086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09966_ (.I(_04086_),
    .Z(_00183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09967_ (.I(_03995_),
    .Z(_04087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09968_ (.A1(_03919_),
    .A2(_04087_),
    .ZN(_04088_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09969_ (.I0(_04073_),
    .I1(\mod.u_cpu.rf_ram.memory[522][0] ),
    .S(_04088_),
    .Z(_04089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09970_ (.I(_04089_),
    .Z(_00184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09971_ (.I(_03762_),
    .Z(_04090_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09972_ (.I(_04090_),
    .Z(_04091_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09973_ (.I0(_04091_),
    .I1(\mod.u_cpu.rf_ram.memory[522][1] ),
    .S(_04088_),
    .Z(_04092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09974_ (.I(_04092_),
    .Z(_00185_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09975_ (.A1(_03714_),
    .A2(_04077_),
    .ZN(_04093_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09976_ (.I0(\mod.u_cpu.rf_ram.memory[521][0] ),
    .I1(_03925_),
    .S(_04093_),
    .Z(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09977_ (.I(_04094_),
    .Z(_00186_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09978_ (.I0(\mod.u_cpu.rf_ram.memory[521][1] ),
    .I1(_03929_),
    .S(_04093_),
    .Z(_04095_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09979_ (.I(_04095_),
    .Z(_00187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09980_ (.I(_04050_),
    .Z(_04096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09981_ (.A1(_03933_),
    .A2(_04087_),
    .ZN(_04097_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09982_ (.I0(_04096_),
    .I1(\mod.u_cpu.rf_ram.memory[520][0] ),
    .S(_04097_),
    .Z(_04098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09983_ (.I(_04098_),
    .Z(_00188_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09984_ (.I0(_04091_),
    .I1(\mod.u_cpu.rf_ram.memory[520][1] ),
    .S(_04097_),
    .Z(_04099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09985_ (.I(_04099_),
    .Z(_00189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09986_ (.A1(_04013_),
    .A2(_03851_),
    .ZN(_04100_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09987_ (.I0(_04096_),
    .I1(\mod.u_cpu.rf_ram.memory[51][0] ),
    .S(_04100_),
    .Z(_04101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09988_ (.I(_04101_),
    .Z(_00190_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09989_ (.I0(_04091_),
    .I1(\mod.u_cpu.rf_ram.memory[51][1] ),
    .S(_04100_),
    .Z(_04102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09990_ (.I(_04102_),
    .Z(_00191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09991_ (.A1(_03951_),
    .A2(_04087_),
    .ZN(_04103_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09992_ (.I0(_04096_),
    .I1(\mod.u_cpu.rf_ram.memory[518][0] ),
    .S(_04103_),
    .Z(_04104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09993_ (.I(_04104_),
    .Z(_00192_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09994_ (.I0(_04091_),
    .I1(\mod.u_cpu.rf_ram.memory[518][1] ),
    .S(_04103_),
    .Z(_04105_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09995_ (.I(_04105_),
    .Z(_00193_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09996_ (.A1(_03702_),
    .A2(_03939_),
    .Z(_04106_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09997_ (.I(_04106_),
    .Z(_04107_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09998_ (.I(_04107_),
    .Z(_04108_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09999_ (.A1(_04077_),
    .A2(_04108_),
    .ZN(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10000_ (.A1(_03899_),
    .A2(_04109_),
    .ZN(_04110_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10001_ (.A1(_02529_),
    .A2(_04109_),
    .B(_04110_),
    .ZN(_00194_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10002_ (.I(_03928_),
    .Z(_04111_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10003_ (.I0(\mod.u_cpu.rf_ram.memory[517][1] ),
    .I1(_04111_),
    .S(_04109_),
    .Z(_04112_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10004_ (.I(_04112_),
    .Z(_00195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10005_ (.A1(_03961_),
    .A2(_04087_),
    .ZN(_04113_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10006_ (.I0(_04096_),
    .I1(\mod.u_cpu.rf_ram.memory[516][0] ),
    .S(_04113_),
    .Z(_04114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10007_ (.I(_04114_),
    .Z(_00196_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10008_ (.I(_04090_),
    .Z(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10009_ (.I0(_04115_),
    .I1(\mod.u_cpu.rf_ram.memory[516][1] ),
    .S(_04113_),
    .Z(_04116_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10010_ (.I(_04116_),
    .Z(_00197_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10011_ (.I(_04050_),
    .Z(_04117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10012_ (.I(_03995_),
    .Z(_04118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10013_ (.A1(_03969_),
    .A2(_04118_),
    .ZN(_04119_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10014_ (.I0(_04117_),
    .I1(\mod.u_cpu.rf_ram.memory[515][0] ),
    .S(_04119_),
    .Z(_04120_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10015_ (.I(_04120_),
    .Z(_00198_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10016_ (.I0(_04115_),
    .I1(\mod.u_cpu.rf_ram.memory[515][1] ),
    .S(_04119_),
    .Z(_04121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10017_ (.I(_04121_),
    .Z(_00199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10018_ (.A1(_03975_),
    .A2(_04118_),
    .ZN(_04122_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10019_ (.I0(_04117_),
    .I1(\mod.u_cpu.rf_ram.memory[514][0] ),
    .S(_04122_),
    .Z(_04123_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10020_ (.I(_04123_),
    .Z(_00200_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10021_ (.I0(_04115_),
    .I1(\mod.u_cpu.rf_ram.memory[514][1] ),
    .S(_04122_),
    .Z(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10022_ (.I(_04124_),
    .Z(_00201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10023_ (.I(_03979_),
    .Z(_04125_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10024_ (.A1(_04125_),
    .A2(_04002_),
    .Z(_04126_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10025_ (.I0(\mod.u_cpu.rf_ram.memory[513][0] ),
    .I1(_03925_),
    .S(_04126_),
    .Z(_04127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10026_ (.I(_04127_),
    .Z(_00202_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10027_ (.I0(\mod.u_cpu.rf_ram.memory[513][1] ),
    .I1(_04111_),
    .S(_04126_),
    .Z(_04128_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10028_ (.I(_04128_),
    .Z(_00203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10029_ (.A1(_03986_),
    .A2(_04118_),
    .ZN(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10030_ (.I0(_04117_),
    .I1(\mod.u_cpu.rf_ram.memory[512][0] ),
    .S(_04129_),
    .Z(_04130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10031_ (.I(_04130_),
    .Z(_00204_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10032_ (.I0(_04115_),
    .I1(\mod.u_cpu.rf_ram.memory[512][1] ),
    .S(_04129_),
    .Z(_04131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10033_ (.I(_04131_),
    .Z(_00205_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10034_ (.A1(_03662_),
    .A2(_03665_),
    .A3(_03753_),
    .ZN(_04132_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10035_ (.A1(\mod.u_cpu.cpu.immdec.imm11_7[2] ),
    .A2(_03715_),
    .A3(_03717_),
    .ZN(_04133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10036_ (.I(_04133_),
    .Z(_04134_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10037_ (.A1(_03992_),
    .A2(_04132_),
    .A3(_04134_),
    .ZN(_04135_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10038_ (.I(_04135_),
    .Z(_04136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10039_ (.I(_04136_),
    .Z(_04137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10040_ (.A1(_03991_),
    .A2(_04137_),
    .ZN(_04138_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10041_ (.A1(_04044_),
    .A2(_04138_),
    .ZN(_04139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10042_ (.A1(_01612_),
    .A2(_04138_),
    .B(_04139_),
    .ZN(_00206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10043_ (.I(_04090_),
    .Z(_04140_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10044_ (.I0(_04140_),
    .I1(\mod.u_cpu.rf_ram.memory[511][1] ),
    .S(_04138_),
    .Z(_04141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10045_ (.I(_04141_),
    .Z(_00207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10046_ (.I(_04135_),
    .Z(_04142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10047_ (.I(_04142_),
    .Z(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10048_ (.A1(_03752_),
    .A2(_04143_),
    .ZN(_04144_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10049_ (.I0(_04117_),
    .I1(\mod.u_cpu.rf_ram.memory[510][0] ),
    .S(_04144_),
    .Z(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10050_ (.I(_04145_),
    .Z(_00208_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10051_ (.I0(_04140_),
    .I1(\mod.u_cpu.rf_ram.memory[510][1] ),
    .S(_04144_),
    .Z(_04146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10052_ (.I(_04146_),
    .Z(_00209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10053_ (.I(_03738_),
    .Z(_04147_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10054_ (.I(_04147_),
    .Z(_04148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10055_ (.A1(_04013_),
    .A2(_03859_),
    .ZN(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10056_ (.I0(_04148_),
    .I1(\mod.u_cpu.rf_ram.memory[50][0] ),
    .S(_04149_),
    .Z(_04150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10057_ (.I(_04150_),
    .Z(_00210_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10058_ (.I0(_04140_),
    .I1(\mod.u_cpu.rf_ram.memory[50][1] ),
    .S(_04149_),
    .Z(_04151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10059_ (.I(_04151_),
    .Z(_00211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10060_ (.A1(_03782_),
    .A2(_04143_),
    .ZN(_04152_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10061_ (.I0(_04148_),
    .I1(\mod.u_cpu.rf_ram.memory[508][0] ),
    .S(_04152_),
    .Z(_04153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10062_ (.I(_04153_),
    .Z(_00212_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10063_ (.I0(_04140_),
    .I1(\mod.u_cpu.rf_ram.memory[508][1] ),
    .S(_04152_),
    .Z(_04154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10064_ (.I(_04154_),
    .Z(_00213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10065_ (.A1(_03791_),
    .A2(_04143_),
    .ZN(_04155_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10066_ (.I0(_04148_),
    .I1(\mod.u_cpu.rf_ram.memory[507][0] ),
    .S(_04155_),
    .Z(_04156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10067_ (.I(_04156_),
    .Z(_00214_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10068_ (.I(_04090_),
    .Z(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10069_ (.I0(_04157_),
    .I1(\mod.u_cpu.rf_ram.memory[507][1] ),
    .S(_04155_),
    .Z(_04158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10070_ (.I(_04158_),
    .Z(_00215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10071_ (.A1(_03797_),
    .A2(_04143_),
    .ZN(_04159_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10072_ (.I0(_04148_),
    .I1(\mod.u_cpu.rf_ram.memory[506][0] ),
    .S(_04159_),
    .Z(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10073_ (.I(_04160_),
    .Z(_00216_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10074_ (.I0(_04157_),
    .I1(\mod.u_cpu.rf_ram.memory[506][1] ),
    .S(_04159_),
    .Z(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10075_ (.I(_04161_),
    .Z(_00217_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10076_ (.I(_04147_),
    .Z(_04162_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10077_ (.I(_04025_),
    .Z(_04163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10078_ (.I(_04142_),
    .Z(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10079_ (.A1(_04163_),
    .A2(_04164_),
    .ZN(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10080_ (.I0(_04162_),
    .I1(\mod.u_cpu.rf_ram.memory[505][0] ),
    .S(_04165_),
    .Z(_04166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10081_ (.I(_04166_),
    .Z(_00218_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10082_ (.I0(_04157_),
    .I1(\mod.u_cpu.rf_ram.memory[505][1] ),
    .S(_04165_),
    .Z(_04167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10083_ (.I(_04167_),
    .Z(_00219_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10084_ (.I(_03804_),
    .Z(_04168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10085_ (.A1(_04168_),
    .A2(_04164_),
    .ZN(_04169_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10086_ (.I0(_04162_),
    .I1(\mod.u_cpu.rf_ram.memory[504][0] ),
    .S(_04169_),
    .Z(_04170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10087_ (.I(_04170_),
    .Z(_00220_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10088_ (.I0(_04157_),
    .I1(\mod.u_cpu.rf_ram.memory[504][1] ),
    .S(_04169_),
    .Z(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10089_ (.I(_04171_),
    .Z(_00221_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10090_ (.I(_03821_),
    .Z(_04172_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10091_ (.I(_04136_),
    .Z(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10092_ (.A1(_04172_),
    .A2(_04173_),
    .ZN(_04174_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10093_ (.A1(_04044_),
    .A2(_04174_),
    .ZN(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10094_ (.A1(_01597_),
    .A2(_04174_),
    .B(_04175_),
    .ZN(_00222_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10095_ (.I(_03761_),
    .Z(_04176_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10096_ (.I(_04176_),
    .Z(_04177_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10097_ (.I(_04177_),
    .Z(_04178_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10098_ (.I0(_04178_),
    .I1(\mod.u_cpu.rf_ram.memory[503][1] ),
    .S(_04174_),
    .Z(_04179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10099_ (.I(_04179_),
    .Z(_00223_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10100_ (.I(_03828_),
    .Z(_04180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10101_ (.A1(_04180_),
    .A2(_04164_),
    .ZN(_04181_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10102_ (.I0(_04162_),
    .I1(\mod.u_cpu.rf_ram.memory[502][0] ),
    .S(_04181_),
    .Z(_04182_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10103_ (.I(_04182_),
    .Z(_00224_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10104_ (.I0(_04178_),
    .I1(\mod.u_cpu.rf_ram.memory[502][1] ),
    .S(_04181_),
    .Z(_04183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10105_ (.I(_04183_),
    .Z(_00225_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10106_ (.I(_03835_),
    .Z(_04184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10107_ (.A1(_04184_),
    .A2(_04173_),
    .ZN(_04185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10108_ (.I(_04043_),
    .Z(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10109_ (.A1(_04186_),
    .A2(_04185_),
    .ZN(_04187_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10110_ (.A1(_01594_),
    .A2(_04185_),
    .B(_04187_),
    .ZN(_00226_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10111_ (.I0(_04178_),
    .I1(\mod.u_cpu.rf_ram.memory[501][1] ),
    .S(_04185_),
    .Z(_04188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10112_ (.I(_04188_),
    .Z(_00227_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10113_ (.I(_03842_),
    .Z(_04189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10114_ (.A1(_04189_),
    .A2(_04164_),
    .ZN(_04190_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10115_ (.I0(_04162_),
    .I1(\mod.u_cpu.rf_ram.memory[500][0] ),
    .S(_04190_),
    .Z(_04191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10116_ (.I(_04191_),
    .Z(_00228_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10117_ (.I0(_04178_),
    .I1(\mod.u_cpu.rf_ram.memory[500][1] ),
    .S(_04190_),
    .Z(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10118_ (.I(_04192_),
    .Z(_00229_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10119_ (.I(_04147_),
    .Z(_04193_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10120_ (.A1(_03722_),
    .A2(_03726_),
    .Z(_04194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10121_ (.I(_04194_),
    .Z(_04195_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10122_ (.I(_04195_),
    .Z(_04196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10123_ (.A1(_04196_),
    .A2(_03961_),
    .ZN(_04197_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10124_ (.I0(_04193_),
    .I1(\mod.u_cpu.rf_ram.memory[4][0] ),
    .S(_04197_),
    .Z(_04198_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10125_ (.I(_04198_),
    .Z(_00230_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10126_ (.I(_04177_),
    .Z(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10127_ (.I0(_04199_),
    .I1(\mod.u_cpu.rf_ram.memory[4][1] ),
    .S(_04197_),
    .Z(_04200_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10128_ (.I(_04200_),
    .Z(_00231_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10129_ (.I(_03858_),
    .Z(_04201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10130_ (.I(_04142_),
    .Z(_04202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10131_ (.A1(_04201_),
    .A2(_04202_),
    .ZN(_04203_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10132_ (.I0(_04193_),
    .I1(\mod.u_cpu.rf_ram.memory[498][0] ),
    .S(_04203_),
    .Z(_04204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10133_ (.I(_04204_),
    .Z(_00232_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10134_ (.I0(_04199_),
    .I1(\mod.u_cpu.rf_ram.memory[498][1] ),
    .S(_04203_),
    .Z(_04205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10135_ (.I(_04205_),
    .Z(_00233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10136_ (.A1(_03866_),
    .A2(_04202_),
    .ZN(_04206_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10137_ (.I0(_04193_),
    .I1(\mod.u_cpu.rf_ram.memory[497][0] ),
    .S(_04206_),
    .Z(_04207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10138_ (.I(_04207_),
    .Z(_00234_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10139_ (.I0(_04199_),
    .I1(\mod.u_cpu.rf_ram.memory[497][1] ),
    .S(_04206_),
    .Z(_04208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10140_ (.I(_04208_),
    .Z(_00235_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10141_ (.I(_03872_),
    .Z(_04209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10142_ (.A1(_04209_),
    .A2(_04202_),
    .ZN(_04210_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10143_ (.I0(_04193_),
    .I1(\mod.u_cpu.rf_ram.memory[496][0] ),
    .S(_04210_),
    .Z(_04211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10144_ (.I(_04211_),
    .Z(_00236_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10145_ (.I0(_04199_),
    .I1(\mod.u_cpu.rf_ram.memory[496][1] ),
    .S(_04210_),
    .Z(_04212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10146_ (.I(_04212_),
    .Z(_00237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10147_ (.A1(_04068_),
    .A2(_04173_),
    .ZN(_04213_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10148_ (.A1(_04186_),
    .A2(_04213_),
    .ZN(_04214_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10149_ (.A1(_01648_),
    .A2(_04213_),
    .B(_04214_),
    .ZN(_00238_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10150_ (.I(_04177_),
    .Z(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10151_ (.I0(_04215_),
    .I1(\mod.u_cpu.rf_ram.memory[495][1] ),
    .S(_04213_),
    .Z(_04216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10152_ (.I(_04216_),
    .Z(_00239_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10153_ (.I(_04147_),
    .Z(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10154_ (.I(_03885_),
    .Z(_04218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10155_ (.A1(_04218_),
    .A2(_04202_),
    .ZN(_04219_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10156_ (.I0(_04217_),
    .I1(\mod.u_cpu.rf_ram.memory[494][0] ),
    .S(_04219_),
    .Z(_04220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10157_ (.I(_04220_),
    .Z(_00240_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10158_ (.I0(_04215_),
    .I1(\mod.u_cpu.rf_ram.memory[494][1] ),
    .S(_04219_),
    .Z(_04221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10159_ (.I(_04221_),
    .Z(_00241_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10160_ (.I(\mod.u_cpu.cpu.immdec.imm11_7[4] ),
    .ZN(_04222_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10161_ (.I(_04222_),
    .Z(_04223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10162_ (.A1(_03662_),
    .A2(_03753_),
    .ZN(_04224_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10163_ (.A1(_04223_),
    .A2(_04224_),
    .ZN(_04225_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10164_ (.A1(_03992_),
    .A2(_04134_),
    .ZN(_04226_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10165_ (.I(_04226_),
    .Z(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10166_ (.A1(_04225_),
    .A2(_04227_),
    .ZN(_04228_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10167_ (.A1(_03896_),
    .A2(_04228_),
    .ZN(_04229_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10168_ (.I(_03898_),
    .Z(_04230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10169_ (.A1(_04230_),
    .A2(_04229_),
    .ZN(_04231_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10170_ (.A1(_01640_),
    .A2(_04229_),
    .B(_04231_),
    .ZN(_00242_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10171_ (.I0(\mod.u_cpu.rf_ram.memory[493][1] ),
    .I1(_04111_),
    .S(_04229_),
    .Z(_04232_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10172_ (.I(_04232_),
    .Z(_00243_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10173_ (.I(_03904_),
    .Z(_04233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10174_ (.I(_04136_),
    .Z(_04234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10175_ (.A1(_04233_),
    .A2(_04234_),
    .ZN(_04235_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10176_ (.I0(_04217_),
    .I1(\mod.u_cpu.rf_ram.memory[492][0] ),
    .S(_04235_),
    .Z(_04236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10177_ (.I(_04236_),
    .Z(_00244_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10178_ (.I0(_04215_),
    .I1(\mod.u_cpu.rf_ram.memory[492][1] ),
    .S(_04235_),
    .Z(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10179_ (.I(_04237_),
    .Z(_00245_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10180_ (.I(_03910_),
    .Z(_04238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10181_ (.A1(_04238_),
    .A2(_04234_),
    .ZN(_04239_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10182_ (.I0(_04217_),
    .I1(\mod.u_cpu.rf_ram.memory[491][0] ),
    .S(_04239_),
    .Z(_04240_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10183_ (.I(_04240_),
    .Z(_00246_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10184_ (.I0(_04215_),
    .I1(\mod.u_cpu.rf_ram.memory[491][1] ),
    .S(_04239_),
    .Z(_04241_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10185_ (.I(_04241_),
    .Z(_00247_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10186_ (.I(_03918_),
    .Z(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10187_ (.A1(_04242_),
    .A2(_04234_),
    .ZN(_04243_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10188_ (.I0(_04217_),
    .I1(\mod.u_cpu.rf_ram.memory[490][0] ),
    .S(_04243_),
    .Z(_04244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10189_ (.I(_04244_),
    .Z(_00248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10190_ (.I(_04177_),
    .Z(_04245_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10191_ (.I0(_04245_),
    .I1(\mod.u_cpu.rf_ram.memory[490][1] ),
    .S(_04243_),
    .Z(_04246_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10192_ (.I(_04246_),
    .Z(_00249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10193_ (.I(_03737_),
    .Z(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10194_ (.I(_04247_),
    .Z(_04248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10195_ (.I(_04248_),
    .Z(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10196_ (.I(_03808_),
    .Z(_04250_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10197_ (.I(_04250_),
    .Z(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10198_ (.A1(_04251_),
    .A2(_03873_),
    .ZN(_04252_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10199_ (.I0(_04249_),
    .I1(\mod.u_cpu.rf_ram.memory[48][0] ),
    .S(_04252_),
    .Z(_04253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10200_ (.I(_04253_),
    .Z(_00250_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10201_ (.I0(_04245_),
    .I1(\mod.u_cpu.rf_ram.memory[48][1] ),
    .S(_04252_),
    .Z(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10202_ (.I(_04254_),
    .Z(_00251_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10203_ (.I(_03932_),
    .Z(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10204_ (.A1(_04255_),
    .A2(_04234_),
    .ZN(_04256_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10205_ (.I0(_04249_),
    .I1(\mod.u_cpu.rf_ram.memory[488][0] ),
    .S(_04256_),
    .Z(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10206_ (.I(_04257_),
    .Z(_00252_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10207_ (.I0(_04245_),
    .I1(\mod.u_cpu.rf_ram.memory[488][1] ),
    .S(_04256_),
    .Z(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10208_ (.I(_04258_),
    .Z(_00253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10209_ (.A1(_03942_),
    .A2(_04173_),
    .ZN(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10210_ (.A1(_04186_),
    .A2(_04259_),
    .ZN(_04260_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10211_ (.A1(_01625_),
    .A2(_04259_),
    .B(_04260_),
    .ZN(_00254_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10212_ (.I0(_04245_),
    .I1(\mod.u_cpu.rf_ram.memory[487][1] ),
    .S(_04259_),
    .Z(_04261_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10213_ (.I(_04261_),
    .Z(_00255_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10214_ (.I(_03950_),
    .Z(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10215_ (.I(_04136_),
    .Z(_04263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10216_ (.A1(_04262_),
    .A2(_04263_),
    .ZN(_04264_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10217_ (.I0(_04249_),
    .I1(\mod.u_cpu.rf_ram.memory[486][0] ),
    .S(_04264_),
    .Z(_04265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10218_ (.I(_04265_),
    .Z(_00256_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10219_ (.I(_04176_),
    .Z(_04266_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10220_ (.I(_04266_),
    .Z(_04267_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10221_ (.I0(_04267_),
    .I1(\mod.u_cpu.rf_ram.memory[486][1] ),
    .S(_04264_),
    .Z(_04268_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10222_ (.I(_04268_),
    .Z(_00257_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10223_ (.A1(_04108_),
    .A2(_04228_),
    .ZN(_04269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10224_ (.A1(_04230_),
    .A2(_04269_),
    .ZN(_04270_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10225_ (.A1(_01622_),
    .A2(_04269_),
    .B(_04270_),
    .ZN(_00258_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10226_ (.I0(\mod.u_cpu.rf_ram.memory[485][1] ),
    .I1(_04111_),
    .S(_04269_),
    .Z(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10227_ (.I(_04271_),
    .Z(_00259_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10228_ (.I(_03960_),
    .Z(_04272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10229_ (.A1(_04272_),
    .A2(_04263_),
    .ZN(_04273_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10230_ (.I0(_04249_),
    .I1(\mod.u_cpu.rf_ram.memory[484][0] ),
    .S(_04273_),
    .Z(_04274_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10231_ (.I(_04274_),
    .Z(_00260_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10232_ (.I0(_04267_),
    .I1(\mod.u_cpu.rf_ram.memory[484][1] ),
    .S(_04273_),
    .Z(_04275_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10233_ (.I(_04275_),
    .Z(_00261_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10234_ (.I(_04248_),
    .Z(_04276_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10235_ (.I(_03968_),
    .Z(_04277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10236_ (.A1(_04277_),
    .A2(_04263_),
    .ZN(_04278_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10237_ (.I0(_04276_),
    .I1(\mod.u_cpu.rf_ram.memory[483][0] ),
    .S(_04278_),
    .Z(_04279_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10238_ (.I(_04279_),
    .Z(_00262_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10239_ (.I0(_04267_),
    .I1(\mod.u_cpu.rf_ram.memory[483][1] ),
    .S(_04278_),
    .Z(_04280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10240_ (.I(_04280_),
    .Z(_00263_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10241_ (.I(_03974_),
    .Z(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10242_ (.A1(_04281_),
    .A2(_04263_),
    .ZN(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10243_ (.I0(_04276_),
    .I1(\mod.u_cpu.rf_ram.memory[482][0] ),
    .S(_04282_),
    .Z(_04283_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10244_ (.I(_04283_),
    .Z(_00264_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10245_ (.I0(_04267_),
    .I1(\mod.u_cpu.rf_ram.memory[482][1] ),
    .S(_04282_),
    .Z(_04284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10246_ (.I(_04284_),
    .Z(_00265_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10247_ (.I(_04125_),
    .Z(_04285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10248_ (.A1(_04285_),
    .A2(_04137_),
    .ZN(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10249_ (.I0(_04276_),
    .I1(\mod.u_cpu.rf_ram.memory[481][0] ),
    .S(_04286_),
    .Z(_04287_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10250_ (.I(_04287_),
    .Z(_00266_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10251_ (.I(_04266_),
    .Z(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10252_ (.I0(_04288_),
    .I1(\mod.u_cpu.rf_ram.memory[481][1] ),
    .S(_04286_),
    .Z(_04289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10253_ (.I(_04289_),
    .Z(_00267_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10254_ (.I(_03985_),
    .Z(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10255_ (.A1(_04290_),
    .A2(_04137_),
    .ZN(_04291_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10256_ (.I0(_04276_),
    .I1(\mod.u_cpu.rf_ram.memory[480][0] ),
    .S(_04291_),
    .Z(_04292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10257_ (.I(_04292_),
    .Z(_00268_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10258_ (.I0(_04288_),
    .I1(\mod.u_cpu.rf_ram.memory[480][1] ),
    .S(_04291_),
    .Z(_04293_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10259_ (.I(_04293_),
    .Z(_00269_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10260_ (.I(_04250_),
    .Z(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10261_ (.A1(_04294_),
    .A2(_04068_),
    .ZN(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10262_ (.A1(_04186_),
    .A2(_04295_),
    .ZN(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10263_ (.A1(_02439_),
    .A2(_04295_),
    .B(_04296_),
    .ZN(_00270_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10264_ (.I0(_04288_),
    .I1(\mod.u_cpu.rf_ram.memory[47][1] ),
    .S(_04295_),
    .Z(_04297_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10265_ (.I(_04297_),
    .Z(_00271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10266_ (.I(_04248_),
    .Z(_04298_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10267_ (.I(_03751_),
    .Z(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10268_ (.A1(_03721_),
    .A2(_04133_),
    .Z(_04300_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10269_ (.A1(_04132_),
    .A2(_04300_),
    .ZN(_04301_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10270_ (.I(_04301_),
    .Z(_04302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10271_ (.I(_04302_),
    .Z(_04303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10272_ (.A1(_04299_),
    .A2(_04303_),
    .ZN(_04304_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10273_ (.I0(_04298_),
    .I1(\mod.u_cpu.rf_ram.memory[478][0] ),
    .S(_04304_),
    .Z(_04305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10274_ (.I(_04305_),
    .Z(_00272_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10275_ (.I0(_04288_),
    .I1(\mod.u_cpu.rf_ram.memory[478][1] ),
    .S(_04304_),
    .Z(_04306_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10276_ (.I(_04306_),
    .Z(_00273_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10277_ (.I(_03769_),
    .Z(_04307_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10278_ (.I(_04301_),
    .Z(_04308_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10279_ (.I(_04308_),
    .Z(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10280_ (.A1(_04307_),
    .A2(_04309_),
    .ZN(_04310_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10281_ (.I(_04043_),
    .Z(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10282_ (.A1(_04311_),
    .A2(_04310_),
    .ZN(_04312_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10283_ (.A1(_01557_),
    .A2(_04310_),
    .B(_04312_),
    .ZN(_00274_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10284_ (.I(_04266_),
    .Z(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10285_ (.I0(_04313_),
    .I1(\mod.u_cpu.rf_ram.memory[477][1] ),
    .S(_04310_),
    .Z(_04314_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10286_ (.I(_04314_),
    .Z(_00275_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10287_ (.I(_03781_),
    .Z(_04315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10288_ (.A1(_04315_),
    .A2(_04303_),
    .ZN(_04316_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10289_ (.I0(_04298_),
    .I1(\mod.u_cpu.rf_ram.memory[476][0] ),
    .S(_04316_),
    .Z(_04317_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10290_ (.I(_04317_),
    .Z(_00276_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10291_ (.I0(_04313_),
    .I1(\mod.u_cpu.rf_ram.memory[476][1] ),
    .S(_04316_),
    .Z(_04318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10292_ (.I(_04318_),
    .Z(_00277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10293_ (.A1(_03791_),
    .A2(_04303_),
    .ZN(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10294_ (.I0(_04298_),
    .I1(\mod.u_cpu.rf_ram.memory[475][0] ),
    .S(_04319_),
    .Z(_04320_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10295_ (.I(_04320_),
    .Z(_00278_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10296_ (.I0(_04313_),
    .I1(\mod.u_cpu.rf_ram.memory[475][1] ),
    .S(_04319_),
    .Z(_04321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10297_ (.I(_04321_),
    .Z(_00279_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10298_ (.I(_03796_),
    .Z(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10299_ (.A1(_04322_),
    .A2(_04303_),
    .ZN(_04323_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10300_ (.I0(_04298_),
    .I1(\mod.u_cpu.rf_ram.memory[474][0] ),
    .S(_04323_),
    .Z(_04324_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10301_ (.I(_04324_),
    .Z(_00280_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10302_ (.I0(_04313_),
    .I1(\mod.u_cpu.rf_ram.memory[474][1] ),
    .S(_04323_),
    .Z(_04325_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10303_ (.I(_04325_),
    .Z(_00281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10304_ (.I(_04248_),
    .Z(_04326_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10305_ (.I(_04302_),
    .Z(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10306_ (.A1(_04163_),
    .A2(_04327_),
    .ZN(_04328_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10307_ (.I0(_04326_),
    .I1(\mod.u_cpu.rf_ram.memory[473][0] ),
    .S(_04328_),
    .Z(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10308_ (.I(_04329_),
    .Z(_00282_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10309_ (.I(_04266_),
    .Z(_04330_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10310_ (.I0(_04330_),
    .I1(\mod.u_cpu.rf_ram.memory[473][1] ),
    .S(_04328_),
    .Z(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10311_ (.I(_04331_),
    .Z(_00283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10312_ (.A1(_04168_),
    .A2(_04327_),
    .ZN(_04332_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10313_ (.I0(_04326_),
    .I1(\mod.u_cpu.rf_ram.memory[472][0] ),
    .S(_04332_),
    .Z(_04333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10314_ (.I(_04333_),
    .Z(_00284_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10315_ (.I0(_04330_),
    .I1(\mod.u_cpu.rf_ram.memory[472][1] ),
    .S(_04332_),
    .Z(_04334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10316_ (.I(_04334_),
    .Z(_00285_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10317_ (.I(_04308_),
    .Z(_04335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10318_ (.A1(_04172_),
    .A2(_04335_),
    .ZN(_04336_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10319_ (.A1(_04311_),
    .A2(_04336_),
    .ZN(_04337_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10320_ (.A1(_01579_),
    .A2(_04336_),
    .B(_04337_),
    .ZN(_00286_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10321_ (.I0(_04330_),
    .I1(\mod.u_cpu.rf_ram.memory[471][1] ),
    .S(_04336_),
    .Z(_04338_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10322_ (.I(_04338_),
    .Z(_00287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10323_ (.A1(_04180_),
    .A2(_04327_),
    .ZN(_04339_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10324_ (.I0(_04326_),
    .I1(\mod.u_cpu.rf_ram.memory[470][0] ),
    .S(_04339_),
    .Z(_04340_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10325_ (.I(_04340_),
    .Z(_00288_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10326_ (.I0(_04330_),
    .I1(\mod.u_cpu.rf_ram.memory[470][1] ),
    .S(_04339_),
    .Z(_04341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10327_ (.I(_04341_),
    .Z(_00289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10328_ (.A1(_04251_),
    .A2(_03886_),
    .ZN(_04342_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10329_ (.I0(_04326_),
    .I1(\mod.u_cpu.rf_ram.memory[46][0] ),
    .S(_04342_),
    .Z(_04343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10330_ (.I(_04343_),
    .Z(_00290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10331_ (.I(_04176_),
    .Z(_04344_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10332_ (.I(_04344_),
    .Z(_04345_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10333_ (.I0(_04345_),
    .I1(\mod.u_cpu.rf_ram.memory[46][1] ),
    .S(_04342_),
    .Z(_04346_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10334_ (.I(_04346_),
    .Z(_00291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10335_ (.I(_04247_),
    .Z(_04347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10336_ (.I(_04347_),
    .Z(_04348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10337_ (.A1(_04189_),
    .A2(_04327_),
    .ZN(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10338_ (.I0(_04348_),
    .I1(\mod.u_cpu.rf_ram.memory[468][0] ),
    .S(_04349_),
    .Z(_04350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10339_ (.I(_04350_),
    .Z(_00292_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10340_ (.I0(_04345_),
    .I1(\mod.u_cpu.rf_ram.memory[468][1] ),
    .S(_04349_),
    .Z(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10341_ (.I(_04351_),
    .Z(_00293_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10342_ (.I(_03850_),
    .Z(_04352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10343_ (.I(_04302_),
    .Z(_04353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10344_ (.A1(_04352_),
    .A2(_04353_),
    .ZN(_04354_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10345_ (.I0(_04348_),
    .I1(\mod.u_cpu.rf_ram.memory[467][0] ),
    .S(_04354_),
    .Z(_04355_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10346_ (.I(_04355_),
    .Z(_00294_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10347_ (.I0(_04345_),
    .I1(\mod.u_cpu.rf_ram.memory[467][1] ),
    .S(_04354_),
    .Z(_04356_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10348_ (.I(_04356_),
    .Z(_00295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10349_ (.A1(_04201_),
    .A2(_04353_),
    .ZN(_04357_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10350_ (.I0(_04348_),
    .I1(\mod.u_cpu.rf_ram.memory[466][0] ),
    .S(_04357_),
    .Z(_04358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10351_ (.I(_04358_),
    .Z(_00296_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10352_ (.I0(_04345_),
    .I1(\mod.u_cpu.rf_ram.memory[466][1] ),
    .S(_04357_),
    .Z(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10353_ (.I(_04359_),
    .Z(_00297_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10354_ (.I(_03865_),
    .Z(_04360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10355_ (.A1(_04360_),
    .A2(_04353_),
    .ZN(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10356_ (.I0(_04348_),
    .I1(\mod.u_cpu.rf_ram.memory[465][0] ),
    .S(_04361_),
    .Z(_04362_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10357_ (.I(_04362_),
    .Z(_00298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10358_ (.I(_04344_),
    .Z(_04363_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10359_ (.I0(_04363_),
    .I1(\mod.u_cpu.rf_ram.memory[465][1] ),
    .S(_04361_),
    .Z(_04364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10360_ (.I(_04364_),
    .Z(_00299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10361_ (.I(_04347_),
    .Z(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10362_ (.A1(_04209_),
    .A2(_04353_),
    .ZN(_04366_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10363_ (.I0(_04365_),
    .I1(\mod.u_cpu.rf_ram.memory[464][0] ),
    .S(_04366_),
    .Z(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10364_ (.I(_04367_),
    .Z(_00300_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10365_ (.I0(_04363_),
    .I1(\mod.u_cpu.rf_ram.memory[464][1] ),
    .S(_04366_),
    .Z(_04368_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10366_ (.I(_04368_),
    .Z(_00301_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10367_ (.I(_04066_),
    .Z(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10368_ (.A1(_04369_),
    .A2(_04335_),
    .ZN(_04370_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10369_ (.A1(_04311_),
    .A2(_04370_),
    .ZN(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10370_ (.A1(_01546_),
    .A2(_04370_),
    .B(_04371_),
    .ZN(_00302_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10371_ (.I0(_04363_),
    .I1(\mod.u_cpu.rf_ram.memory[463][1] ),
    .S(_04370_),
    .Z(_04372_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10372_ (.I(_04372_),
    .Z(_00303_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10373_ (.I(_04308_),
    .Z(_04373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10374_ (.A1(_04218_),
    .A2(_04373_),
    .ZN(_04374_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10375_ (.I0(_04365_),
    .I1(\mod.u_cpu.rf_ram.memory[462][0] ),
    .S(_04374_),
    .Z(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10376_ (.I(_04375_),
    .Z(_00304_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10377_ (.I0(_04363_),
    .I1(\mod.u_cpu.rf_ram.memory[462][1] ),
    .S(_04374_),
    .Z(_04376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10378_ (.I(_04376_),
    .Z(_00305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10379_ (.I(_03894_),
    .Z(_04377_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10380_ (.A1(_03721_),
    .A2(_04134_),
    .ZN(_04378_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10381_ (.I(_04378_),
    .Z(_04379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10382_ (.A1(_04225_),
    .A2(_04379_),
    .ZN(_04380_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10383_ (.A1(_04377_),
    .A2(_04380_),
    .ZN(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10384_ (.A1(_04230_),
    .A2(_04381_),
    .ZN(_04382_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10385_ (.A1(_01542_),
    .A2(_04381_),
    .B(_04382_),
    .ZN(_00306_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10386_ (.I(_03928_),
    .Z(_04383_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10387_ (.I0(\mod.u_cpu.rf_ram.memory[461][1] ),
    .I1(_04383_),
    .S(_04381_),
    .Z(_04384_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10388_ (.I(_04384_),
    .Z(_00307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10389_ (.A1(_04233_),
    .A2(_04373_),
    .ZN(_04385_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10390_ (.I0(_04365_),
    .I1(\mod.u_cpu.rf_ram.memory[460][0] ),
    .S(_04385_),
    .Z(_04386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10391_ (.I(_04386_),
    .Z(_00308_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10392_ (.I(_04344_),
    .Z(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10393_ (.I0(_04387_),
    .I1(\mod.u_cpu.rf_ram.memory[460][1] ),
    .S(_04385_),
    .Z(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10394_ (.I(_04388_),
    .Z(_00309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10395_ (.A1(_03727_),
    .A2(_03807_),
    .ZN(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10396_ (.A1(_04389_),
    .A2(_03896_),
    .ZN(_04390_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10397_ (.A1(_04230_),
    .A2(_04390_),
    .ZN(_04391_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10398_ (.A1(_02436_),
    .A2(_04390_),
    .B(_04391_),
    .ZN(_00310_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10399_ (.I0(\mod.u_cpu.rf_ram.memory[45][1] ),
    .I1(_04383_),
    .S(_04390_),
    .Z(_04392_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10400_ (.I(_04392_),
    .Z(_00311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10401_ (.A1(_04242_),
    .A2(_04373_),
    .ZN(_04393_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10402_ (.I0(_04365_),
    .I1(\mod.u_cpu.rf_ram.memory[458][0] ),
    .S(_04393_),
    .Z(_04394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10403_ (.I(_04394_),
    .Z(_00312_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10404_ (.I0(_04387_),
    .I1(\mod.u_cpu.rf_ram.memory[458][1] ),
    .S(_04393_),
    .Z(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10405_ (.I(_04395_),
    .Z(_00313_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10406_ (.I(_03924_),
    .Z(_04396_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10407_ (.A1(_03714_),
    .A2(_04380_),
    .ZN(_04397_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10408_ (.I0(\mod.u_cpu.rf_ram.memory[457][0] ),
    .I1(_04396_),
    .S(_04397_),
    .Z(_04398_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10409_ (.I(_04398_),
    .Z(_00314_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10410_ (.I0(\mod.u_cpu.rf_ram.memory[457][1] ),
    .I1(_04383_),
    .S(_04397_),
    .Z(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10411_ (.I(_04399_),
    .Z(_00315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10412_ (.I(_04347_),
    .Z(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10413_ (.A1(_04255_),
    .A2(_04373_),
    .ZN(_04401_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10414_ (.I0(_04400_),
    .I1(\mod.u_cpu.rf_ram.memory[456][0] ),
    .S(_04401_),
    .Z(_04402_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10415_ (.I(_04402_),
    .Z(_00316_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10416_ (.I0(_04387_),
    .I1(\mod.u_cpu.rf_ram.memory[456][1] ),
    .S(_04401_),
    .Z(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10417_ (.I(_04403_),
    .Z(_00317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10418_ (.A1(_03942_),
    .A2(_04335_),
    .ZN(_04404_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10419_ (.A1(_04311_),
    .A2(_04404_),
    .ZN(_04405_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10420_ (.A1(_01521_),
    .A2(_04404_),
    .B(_04405_),
    .ZN(_00318_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10421_ (.I0(_04387_),
    .I1(\mod.u_cpu.rf_ram.memory[455][1] ),
    .S(_04404_),
    .Z(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10422_ (.I(_04406_),
    .Z(_00319_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10423_ (.I(_04308_),
    .Z(_04407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10424_ (.A1(_04262_),
    .A2(_04407_),
    .ZN(_04408_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10425_ (.I0(_04400_),
    .I1(\mod.u_cpu.rf_ram.memory[454][0] ),
    .S(_04408_),
    .Z(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10426_ (.I(_04409_),
    .Z(_00320_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10427_ (.I(_04344_),
    .Z(_04410_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10428_ (.I0(_04410_),
    .I1(\mod.u_cpu.rf_ram.memory[454][1] ),
    .S(_04408_),
    .Z(_04411_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10429_ (.I(_04411_),
    .Z(_00321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10430_ (.I(_04106_),
    .Z(_04412_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10431_ (.A1(_04412_),
    .A2(_04380_),
    .ZN(_04413_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10432_ (.I(_03898_),
    .Z(_04414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10433_ (.A1(_04414_),
    .A2(_04413_),
    .ZN(_04415_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10434_ (.A1(_01512_),
    .A2(_04413_),
    .B(_04415_),
    .ZN(_00322_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10435_ (.I0(\mod.u_cpu.rf_ram.memory[453][1] ),
    .I1(_04383_),
    .S(_04413_),
    .Z(_04416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10436_ (.I(_04416_),
    .Z(_00323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10437_ (.A1(_04272_),
    .A2(_04407_),
    .ZN(_04417_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10438_ (.I0(_04400_),
    .I1(\mod.u_cpu.rf_ram.memory[452][0] ),
    .S(_04417_),
    .Z(_04418_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10439_ (.I(_04418_),
    .Z(_00324_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10440_ (.I0(_04410_),
    .I1(\mod.u_cpu.rf_ram.memory[452][1] ),
    .S(_04417_),
    .Z(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10441_ (.I(_04419_),
    .Z(_00325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10442_ (.A1(_04277_),
    .A2(_04407_),
    .ZN(_04420_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10443_ (.I0(_04400_),
    .I1(\mod.u_cpu.rf_ram.memory[451][0] ),
    .S(_04420_),
    .Z(_04421_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10444_ (.I(_04421_),
    .Z(_00326_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10445_ (.I0(_04410_),
    .I1(\mod.u_cpu.rf_ram.memory[451][1] ),
    .S(_04420_),
    .Z(_04422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10446_ (.I(_04422_),
    .Z(_00327_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10447_ (.I(_04347_),
    .Z(_04423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10448_ (.A1(_04281_),
    .A2(_04407_),
    .ZN(_04424_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10449_ (.I0(_04423_),
    .I1(\mod.u_cpu.rf_ram.memory[450][0] ),
    .S(_04424_),
    .Z(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10450_ (.I(_04425_),
    .Z(_00328_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10451_ (.I0(_04410_),
    .I1(\mod.u_cpu.rf_ram.memory[450][1] ),
    .S(_04424_),
    .Z(_04426_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10452_ (.I(_04426_),
    .Z(_00329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10453_ (.A1(_04251_),
    .A2(_03905_),
    .ZN(_04427_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10454_ (.I0(_04423_),
    .I1(\mod.u_cpu.rf_ram.memory[44][0] ),
    .S(_04427_),
    .Z(_04428_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10455_ (.I(_04428_),
    .Z(_00330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10456_ (.I(_04176_),
    .Z(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10457_ (.I(_04429_),
    .Z(_04430_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10458_ (.I0(_04430_),
    .I1(\mod.u_cpu.rf_ram.memory[44][1] ),
    .S(_04427_),
    .Z(_04431_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10459_ (.I(_04431_),
    .Z(_00331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10460_ (.A1(_04290_),
    .A2(_04309_),
    .ZN(_04432_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10461_ (.I0(_04423_),
    .I1(\mod.u_cpu.rf_ram.memory[448][0] ),
    .S(_04432_),
    .Z(_04433_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10462_ (.I(_04433_),
    .Z(_00332_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10463_ (.I0(_04430_),
    .I1(\mod.u_cpu.rf_ram.memory[448][1] ),
    .S(_04432_),
    .Z(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10464_ (.I(_04434_),
    .Z(_00333_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10465_ (.A1(_03755_),
    .A2(_04132_),
    .ZN(_04435_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10466_ (.I(_04435_),
    .Z(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10467_ (.I(_04436_),
    .Z(_04437_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10468_ (.A1(_03991_),
    .A2(_04437_),
    .ZN(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10469_ (.I(_04043_),
    .Z(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10470_ (.A1(_04439_),
    .A2(_04438_),
    .ZN(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10471_ (.A1(_01808_),
    .A2(_04438_),
    .B(_04440_),
    .ZN(_00334_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10472_ (.I0(_04430_),
    .I1(\mod.u_cpu.rf_ram.memory[447][1] ),
    .S(_04438_),
    .Z(_04441_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10473_ (.I(_04441_),
    .Z(_00335_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10474_ (.I(_04435_),
    .Z(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10475_ (.I(_04442_),
    .Z(_04443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10476_ (.A1(_04299_),
    .A2(_04443_),
    .ZN(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10477_ (.I0(_04423_),
    .I1(\mod.u_cpu.rf_ram.memory[446][0] ),
    .S(_04444_),
    .Z(_04445_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10478_ (.I(_04445_),
    .Z(_00336_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10479_ (.I0(_04430_),
    .I1(\mod.u_cpu.rf_ram.memory[446][1] ),
    .S(_04444_),
    .Z(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10480_ (.I(_04446_),
    .Z(_00337_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10481_ (.I(_04436_),
    .Z(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10482_ (.A1(_04307_),
    .A2(_04447_),
    .ZN(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10483_ (.A1(_04439_),
    .A2(_04448_),
    .ZN(_04449_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10484_ (.A1(_01803_),
    .A2(_04448_),
    .B(_04449_),
    .ZN(_00338_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10485_ (.I(_04429_),
    .Z(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10486_ (.I0(_04450_),
    .I1(\mod.u_cpu.rf_ram.memory[445][1] ),
    .S(_04448_),
    .Z(_04451_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10487_ (.I(_04451_),
    .Z(_00339_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10488_ (.I(_04247_),
    .Z(_04452_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10489_ (.I(_04452_),
    .Z(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10490_ (.A1(_04315_),
    .A2(_04443_),
    .ZN(_04454_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10491_ (.I0(_04453_),
    .I1(\mod.u_cpu.rf_ram.memory[444][0] ),
    .S(_04454_),
    .Z(_04455_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10492_ (.I(_04455_),
    .Z(_00340_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10493_ (.I0(_04450_),
    .I1(\mod.u_cpu.rf_ram.memory[444][1] ),
    .S(_04454_),
    .Z(_04456_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10494_ (.I(_04456_),
    .Z(_00341_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10495_ (.I(_03790_),
    .Z(_04457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10496_ (.A1(_04457_),
    .A2(_04443_),
    .ZN(_04458_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10497_ (.I0(_04453_),
    .I1(\mod.u_cpu.rf_ram.memory[443][0] ),
    .S(_04458_),
    .Z(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10498_ (.I(_04459_),
    .Z(_00342_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10499_ (.I0(_04450_),
    .I1(\mod.u_cpu.rf_ram.memory[443][1] ),
    .S(_04458_),
    .Z(_04460_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10500_ (.I(_04460_),
    .Z(_00343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10501_ (.A1(_04322_),
    .A2(_04443_),
    .ZN(_04461_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10502_ (.I0(_04453_),
    .I1(\mod.u_cpu.rf_ram.memory[442][0] ),
    .S(_04461_),
    .Z(_04462_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10503_ (.I(_04462_),
    .Z(_00344_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10504_ (.I0(_04450_),
    .I1(\mod.u_cpu.rf_ram.memory[442][1] ),
    .S(_04461_),
    .Z(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10505_ (.I(_04463_),
    .Z(_00345_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10506_ (.I(_04442_),
    .Z(_04464_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10507_ (.A1(_04163_),
    .A2(_04464_),
    .ZN(_04465_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10508_ (.I0(_04453_),
    .I1(\mod.u_cpu.rf_ram.memory[441][0] ),
    .S(_04465_),
    .Z(_04466_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10509_ (.I(_04466_),
    .Z(_00346_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10510_ (.I(_04429_),
    .Z(_04467_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10511_ (.I0(_04467_),
    .I1(\mod.u_cpu.rf_ram.memory[441][1] ),
    .S(_04465_),
    .Z(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10512_ (.I(_04468_),
    .Z(_00347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10513_ (.I(_04452_),
    .Z(_04469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10514_ (.A1(_04168_),
    .A2(_04464_),
    .ZN(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10515_ (.I0(_04469_),
    .I1(\mod.u_cpu.rf_ram.memory[440][0] ),
    .S(_04470_),
    .Z(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10516_ (.I(_04471_),
    .Z(_00348_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10517_ (.I0(_04467_),
    .I1(\mod.u_cpu.rf_ram.memory[440][1] ),
    .S(_04470_),
    .Z(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10518_ (.I(_04472_),
    .Z(_00349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10519_ (.A1(_04251_),
    .A2(_03911_),
    .ZN(_04473_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10520_ (.I0(_04469_),
    .I1(\mod.u_cpu.rf_ram.memory[43][0] ),
    .S(_04473_),
    .Z(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10521_ (.I(_04474_),
    .Z(_00350_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10522_ (.I0(_04467_),
    .I1(\mod.u_cpu.rf_ram.memory[43][1] ),
    .S(_04473_),
    .Z(_04475_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10523_ (.I(_04475_),
    .Z(_00351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10524_ (.A1(_04180_),
    .A2(_04464_),
    .ZN(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10525_ (.I0(_04469_),
    .I1(\mod.u_cpu.rf_ram.memory[438][0] ),
    .S(_04476_),
    .Z(_04477_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10526_ (.I(_04477_),
    .Z(_00352_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10527_ (.I0(_04467_),
    .I1(\mod.u_cpu.rf_ram.memory[438][1] ),
    .S(_04476_),
    .Z(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10528_ (.I(_04478_),
    .Z(_00353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10529_ (.A1(_04184_),
    .A2(_04447_),
    .ZN(_04479_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10530_ (.A1(_04439_),
    .A2(_04479_),
    .ZN(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10531_ (.A1(_01793_),
    .A2(_04479_),
    .B(_04480_),
    .ZN(_00354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10532_ (.I(_04429_),
    .Z(_04481_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10533_ (.I0(_04481_),
    .I1(\mod.u_cpu.rf_ram.memory[437][1] ),
    .S(_04479_),
    .Z(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10534_ (.I(_04482_),
    .Z(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10535_ (.A1(_04189_),
    .A2(_04464_),
    .ZN(_04483_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10536_ (.I0(_04469_),
    .I1(\mod.u_cpu.rf_ram.memory[436][0] ),
    .S(_04483_),
    .Z(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10537_ (.I(_04484_),
    .Z(_00356_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10538_ (.I0(_04481_),
    .I1(\mod.u_cpu.rf_ram.memory[436][1] ),
    .S(_04483_),
    .Z(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10539_ (.I(_04485_),
    .Z(_00357_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10540_ (.I(_04452_),
    .Z(_04486_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10541_ (.I(_04442_),
    .Z(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10542_ (.A1(_04352_),
    .A2(_04487_),
    .ZN(_04488_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10543_ (.I0(_04486_),
    .I1(\mod.u_cpu.rf_ram.memory[435][0] ),
    .S(_04488_),
    .Z(_04489_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10544_ (.I(_04489_),
    .Z(_00358_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10545_ (.I0(_04481_),
    .I1(\mod.u_cpu.rf_ram.memory[435][1] ),
    .S(_04488_),
    .Z(_04490_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10546_ (.I(_04490_),
    .Z(_00359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10547_ (.A1(_04201_),
    .A2(_04487_),
    .ZN(_04491_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10548_ (.I0(_04486_),
    .I1(\mod.u_cpu.rf_ram.memory[434][0] ),
    .S(_04491_),
    .Z(_04492_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10549_ (.I(_04492_),
    .Z(_00360_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10550_ (.I0(_04481_),
    .I1(\mod.u_cpu.rf_ram.memory[434][1] ),
    .S(_04491_),
    .Z(_04493_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10551_ (.I(_04493_),
    .Z(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10552_ (.A1(_04360_),
    .A2(_04487_),
    .ZN(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10553_ (.I0(_04486_),
    .I1(\mod.u_cpu.rf_ram.memory[433][0] ),
    .S(_04494_),
    .Z(_04495_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10554_ (.I(_04495_),
    .Z(_00362_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10555_ (.I(_03761_),
    .Z(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10556_ (.I(_04496_),
    .Z(_04497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10557_ (.I(_04497_),
    .Z(_04498_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10558_ (.I0(_04498_),
    .I1(\mod.u_cpu.rf_ram.memory[433][1] ),
    .S(_04494_),
    .Z(_04499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10559_ (.I(_04499_),
    .Z(_00363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10560_ (.A1(_04209_),
    .A2(_04487_),
    .ZN(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10561_ (.I0(_04486_),
    .I1(\mod.u_cpu.rf_ram.memory[432][0] ),
    .S(_04500_),
    .Z(_04501_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10562_ (.I(_04501_),
    .Z(_00364_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10563_ (.I0(_04498_),
    .I1(\mod.u_cpu.rf_ram.memory[432][1] ),
    .S(_04500_),
    .Z(_04502_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10564_ (.I(_04502_),
    .Z(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10565_ (.A1(_04369_),
    .A2(_04447_),
    .ZN(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10566_ (.A1(_04439_),
    .A2(_04503_),
    .ZN(_04504_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10567_ (.A1(_01780_),
    .A2(_04503_),
    .B(_04504_),
    .ZN(_00366_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10568_ (.I0(_04498_),
    .I1(\mod.u_cpu.rf_ram.memory[431][1] ),
    .S(_04503_),
    .Z(_04505_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10569_ (.I(_04505_),
    .Z(_00367_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10570_ (.I(_04452_),
    .Z(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10571_ (.I(_04436_),
    .Z(_04507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10572_ (.A1(_04218_),
    .A2(_04507_),
    .ZN(_04508_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10573_ (.I0(_04506_),
    .I1(\mod.u_cpu.rf_ram.memory[430][0] ),
    .S(_04508_),
    .Z(_04509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10574_ (.I(_04509_),
    .Z(_00368_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10575_ (.I0(_04498_),
    .I1(\mod.u_cpu.rf_ram.memory[430][1] ),
    .S(_04508_),
    .Z(_04510_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10576_ (.I(_04510_),
    .Z(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10577_ (.I(_04250_),
    .Z(_04511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10578_ (.A1(_04511_),
    .A2(_03919_),
    .ZN(_04512_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10579_ (.I0(_04506_),
    .I1(\mod.u_cpu.rf_ram.memory[42][0] ),
    .S(_04512_),
    .Z(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10580_ (.I(_04513_),
    .Z(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10581_ (.I(_04497_),
    .Z(_04514_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10582_ (.I0(_04514_),
    .I1(\mod.u_cpu.rf_ram.memory[42][1] ),
    .S(_04512_),
    .Z(_04515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10583_ (.I(_04515_),
    .Z(_00371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10584_ (.A1(_04233_),
    .A2(_04507_),
    .ZN(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10585_ (.I0(_04506_),
    .I1(\mod.u_cpu.rf_ram.memory[428][0] ),
    .S(_04516_),
    .Z(_04517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10586_ (.I(_04517_),
    .Z(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10587_ (.I0(_04514_),
    .I1(\mod.u_cpu.rf_ram.memory[428][1] ),
    .S(_04516_),
    .Z(_04518_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10588_ (.I(_04518_),
    .Z(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10589_ (.A1(_04238_),
    .A2(_04507_),
    .ZN(_04519_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10590_ (.I0(_04506_),
    .I1(\mod.u_cpu.rf_ram.memory[427][0] ),
    .S(_04519_),
    .Z(_04520_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10591_ (.I(_04520_),
    .Z(_00374_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10592_ (.I0(_04514_),
    .I1(\mod.u_cpu.rf_ram.memory[427][1] ),
    .S(_04519_),
    .Z(_04521_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10593_ (.I(_04521_),
    .Z(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10594_ (.I(_04247_),
    .Z(_04522_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10595_ (.I(_04522_),
    .Z(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10596_ (.A1(_04242_),
    .A2(_04507_),
    .ZN(_04524_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10597_ (.I0(_04523_),
    .I1(\mod.u_cpu.rf_ram.memory[426][0] ),
    .S(_04524_),
    .Z(_04525_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10598_ (.I(_04525_),
    .Z(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10599_ (.I0(_04514_),
    .I1(\mod.u_cpu.rf_ram.memory[426][1] ),
    .S(_04524_),
    .Z(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10600_ (.I(_04526_),
    .Z(_00377_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10601_ (.I(_03713_),
    .Z(_04527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10602_ (.A1(_03892_),
    .A2(_04225_),
    .ZN(_04528_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10603_ (.A1(_04527_),
    .A2(_04528_),
    .ZN(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10604_ (.I0(\mod.u_cpu.rf_ram.memory[425][0] ),
    .I1(_04396_),
    .S(_04529_),
    .Z(_04530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10605_ (.I(_04530_),
    .Z(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10606_ (.I(_03733_),
    .Z(_04531_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10607_ (.I(_04531_),
    .Z(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10608_ (.I0(\mod.u_cpu.rf_ram.memory[425][1] ),
    .I1(_04532_),
    .S(_04529_),
    .Z(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10609_ (.I(_04533_),
    .Z(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10610_ (.I(_04436_),
    .Z(_04534_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10611_ (.A1(_04255_),
    .A2(_04534_),
    .ZN(_04535_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10612_ (.I0(_04523_),
    .I1(\mod.u_cpu.rf_ram.memory[424][0] ),
    .S(_04535_),
    .Z(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10613_ (.I(_04536_),
    .Z(_00380_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10614_ (.I(_04497_),
    .Z(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10615_ (.I0(_04537_),
    .I1(\mod.u_cpu.rf_ram.memory[424][1] ),
    .S(_04535_),
    .Z(_04538_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10616_ (.I(_04538_),
    .Z(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10617_ (.I(_03940_),
    .Z(_04539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10618_ (.A1(_04539_),
    .A2(_04447_),
    .ZN(_04540_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10619_ (.I(_03773_),
    .Z(_04541_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10620_ (.I(_04541_),
    .Z(_04542_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10621_ (.A1(_04542_),
    .A2(_04540_),
    .ZN(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10622_ (.A1(_01760_),
    .A2(_04540_),
    .B(_04543_),
    .ZN(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10623_ (.I0(_04537_),
    .I1(\mod.u_cpu.rf_ram.memory[423][1] ),
    .S(_04540_),
    .Z(_04544_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10624_ (.I(_04544_),
    .Z(_00383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10625_ (.A1(_04262_),
    .A2(_04534_),
    .ZN(_04545_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10626_ (.I0(_04523_),
    .I1(\mod.u_cpu.rf_ram.memory[422][0] ),
    .S(_04545_),
    .Z(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10627_ (.I(_04546_),
    .Z(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10628_ (.I0(_04537_),
    .I1(\mod.u_cpu.rf_ram.memory[422][1] ),
    .S(_04545_),
    .Z(_04547_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10629_ (.I(_04547_),
    .Z(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10630_ (.A1(_04412_),
    .A2(_04528_),
    .ZN(_04548_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10631_ (.A1(_04414_),
    .A2(_04548_),
    .ZN(_04549_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10632_ (.A1(_01754_),
    .A2(_04548_),
    .B(_04549_),
    .ZN(_00386_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10633_ (.I0(\mod.u_cpu.rf_ram.memory[421][1] ),
    .I1(_04532_),
    .S(_04548_),
    .Z(_04550_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10634_ (.I(_04550_),
    .Z(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10635_ (.A1(_04272_),
    .A2(_04534_),
    .ZN(_04551_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10636_ (.I0(_04523_),
    .I1(\mod.u_cpu.rf_ram.memory[420][0] ),
    .S(_04551_),
    .Z(_04552_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10637_ (.I(_04552_),
    .Z(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10638_ (.I0(_04537_),
    .I1(\mod.u_cpu.rf_ram.memory[420][1] ),
    .S(_04551_),
    .Z(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10639_ (.I(_04553_),
    .Z(_00389_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10640_ (.A1(_04527_),
    .A2(_04389_),
    .ZN(_04554_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10641_ (.I0(\mod.u_cpu.rf_ram.memory[41][0] ),
    .I1(_04396_),
    .S(_04554_),
    .Z(_04555_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10642_ (.I(_04555_),
    .Z(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10643_ (.I0(\mod.u_cpu.rf_ram.memory[41][1] ),
    .I1(_04532_),
    .S(_04554_),
    .Z(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10644_ (.I(_04556_),
    .Z(_00391_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10645_ (.I(_04522_),
    .Z(_04557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10646_ (.A1(_04281_),
    .A2(_04534_),
    .ZN(_04558_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10647_ (.I0(_04557_),
    .I1(\mod.u_cpu.rf_ram.memory[418][0] ),
    .S(_04558_),
    .Z(_04559_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10648_ (.I(_04559_),
    .Z(_00392_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10649_ (.I(_04497_),
    .Z(_04560_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10650_ (.I0(_04560_),
    .I1(\mod.u_cpu.rf_ram.memory[418][1] ),
    .S(_04558_),
    .Z(_04561_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10651_ (.I(_04561_),
    .Z(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10652_ (.A1(_04285_),
    .A2(_04437_),
    .ZN(_04562_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10653_ (.I0(_04557_),
    .I1(\mod.u_cpu.rf_ram.memory[417][0] ),
    .S(_04562_),
    .Z(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10654_ (.I(_04563_),
    .Z(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10655_ (.I0(_04560_),
    .I1(\mod.u_cpu.rf_ram.memory[417][1] ),
    .S(_04562_),
    .Z(_04564_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10656_ (.I(_04564_),
    .Z(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10657_ (.A1(_04290_),
    .A2(_04437_),
    .ZN(_04565_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10658_ (.I0(_04557_),
    .I1(\mod.u_cpu.rf_ram.memory[416][0] ),
    .S(_04565_),
    .Z(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10659_ (.I(_04566_),
    .Z(_00396_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10660_ (.I0(_04560_),
    .I1(\mod.u_cpu.rf_ram.memory[416][1] ),
    .S(_04565_),
    .Z(_04567_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10661_ (.I(_04567_),
    .Z(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10662_ (.A1(_03993_),
    .A2(_04132_),
    .ZN(_04568_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10663_ (.I(_04568_),
    .Z(_04569_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10664_ (.I(_04569_),
    .Z(_04570_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10665_ (.A1(_03991_),
    .A2(_04570_),
    .ZN(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10666_ (.A1(_04542_),
    .A2(_04571_),
    .ZN(_04572_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10667_ (.A1(_01712_),
    .A2(_04571_),
    .B(_04572_),
    .ZN(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10668_ (.I0(_04560_),
    .I1(\mod.u_cpu.rf_ram.memory[415][1] ),
    .S(_04571_),
    .Z(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10669_ (.I(_04573_),
    .Z(_00399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10670_ (.I(_04568_),
    .Z(_04574_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10671_ (.I(_04574_),
    .Z(_04575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10672_ (.A1(_04299_),
    .A2(_04575_),
    .ZN(_04576_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10673_ (.I0(_04557_),
    .I1(\mod.u_cpu.rf_ram.memory[414][0] ),
    .S(_04576_),
    .Z(_04577_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10674_ (.I(_04577_),
    .Z(_00400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10675_ (.I(_04496_),
    .Z(_04578_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10676_ (.I(_04578_),
    .Z(_04579_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10677_ (.I0(_04579_),
    .I1(\mod.u_cpu.rf_ram.memory[414][1] ),
    .S(_04576_),
    .Z(_04580_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10678_ (.I(_04580_),
    .Z(_00401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10679_ (.A1(_04307_),
    .A2(_04570_),
    .ZN(_04581_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10680_ (.A1(_04542_),
    .A2(_04581_),
    .ZN(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10681_ (.A1(_01706_),
    .A2(_04581_),
    .B(_04582_),
    .ZN(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10682_ (.I0(_04579_),
    .I1(\mod.u_cpu.rf_ram.memory[413][1] ),
    .S(_04581_),
    .Z(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10683_ (.I(_04583_),
    .Z(_00403_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10684_ (.I(_04522_),
    .Z(_04584_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10685_ (.A1(_04315_),
    .A2(_04575_),
    .ZN(_04585_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10686_ (.I0(_04584_),
    .I1(\mod.u_cpu.rf_ram.memory[412][0] ),
    .S(_04585_),
    .Z(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10687_ (.I(_04586_),
    .Z(_00404_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10688_ (.I0(_04579_),
    .I1(\mod.u_cpu.rf_ram.memory[412][1] ),
    .S(_04585_),
    .Z(_04587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10689_ (.I(_04587_),
    .Z(_00405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10690_ (.A1(_04457_),
    .A2(_04575_),
    .ZN(_04588_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10691_ (.I0(_04584_),
    .I1(\mod.u_cpu.rf_ram.memory[411][0] ),
    .S(_04588_),
    .Z(_04589_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10692_ (.I(_04589_),
    .Z(_00406_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10693_ (.I0(_04579_),
    .I1(\mod.u_cpu.rf_ram.memory[411][1] ),
    .S(_04588_),
    .Z(_04590_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10694_ (.I(_04590_),
    .Z(_00407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10695_ (.A1(_04322_),
    .A2(_04575_),
    .ZN(_04591_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10696_ (.I0(_04584_),
    .I1(\mod.u_cpu.rf_ram.memory[410][0] ),
    .S(_04591_),
    .Z(_04592_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10697_ (.I(_04592_),
    .Z(_00408_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10698_ (.I(_04578_),
    .Z(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10699_ (.I0(_04593_),
    .I1(\mod.u_cpu.rf_ram.memory[410][1] ),
    .S(_04591_),
    .Z(_04594_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10700_ (.I(_04594_),
    .Z(_00409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10701_ (.A1(_04511_),
    .A2(_03933_),
    .ZN(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10702_ (.I0(_04584_),
    .I1(\mod.u_cpu.rf_ram.memory[40][0] ),
    .S(_04595_),
    .Z(_04596_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10703_ (.I(_04596_),
    .Z(_00410_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10704_ (.I0(_04593_),
    .I1(\mod.u_cpu.rf_ram.memory[40][1] ),
    .S(_04595_),
    .Z(_04597_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10705_ (.I(_04597_),
    .Z(_00411_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10706_ (.I(_04522_),
    .Z(_04598_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10707_ (.I(_04574_),
    .Z(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10708_ (.A1(_04168_),
    .A2(_04599_),
    .ZN(_04600_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10709_ (.I0(_04598_),
    .I1(\mod.u_cpu.rf_ram.memory[408][0] ),
    .S(_04600_),
    .Z(_04601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10710_ (.I(_04601_),
    .Z(_00412_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10711_ (.I0(_04593_),
    .I1(\mod.u_cpu.rf_ram.memory[408][1] ),
    .S(_04600_),
    .Z(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10712_ (.I(_04602_),
    .Z(_00413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10713_ (.A1(_04172_),
    .A2(_04570_),
    .ZN(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10714_ (.A1(_04542_),
    .A2(_04603_),
    .ZN(_04604_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10715_ (.A1(_01730_),
    .A2(_04603_),
    .B(_04604_),
    .ZN(_00414_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10716_ (.I0(_04593_),
    .I1(\mod.u_cpu.rf_ram.memory[407][1] ),
    .S(_04603_),
    .Z(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10717_ (.I(_04605_),
    .Z(_00415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10718_ (.A1(_04180_),
    .A2(_04599_),
    .ZN(_04606_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10719_ (.I0(_04598_),
    .I1(\mod.u_cpu.rf_ram.memory[406][0] ),
    .S(_04606_),
    .Z(_04607_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10720_ (.I(_04607_),
    .Z(_00416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10721_ (.I(_04578_),
    .Z(_04608_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10722_ (.I0(_04608_),
    .I1(\mod.u_cpu.rf_ram.memory[406][1] ),
    .S(_04606_),
    .Z(_04609_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10723_ (.I(_04609_),
    .Z(_00417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10724_ (.A1(_04184_),
    .A2(_04574_),
    .ZN(_04610_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10725_ (.I(_04541_),
    .Z(_04611_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10726_ (.A1(_04611_),
    .A2(_04610_),
    .ZN(_04612_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10727_ (.A1(_01725_),
    .A2(_04610_),
    .B(_04612_),
    .ZN(_00418_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10728_ (.I0(_04608_),
    .I1(\mod.u_cpu.rf_ram.memory[405][1] ),
    .S(_04610_),
    .Z(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10729_ (.I(_04613_),
    .Z(_00419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10730_ (.A1(_04189_),
    .A2(_04599_),
    .ZN(_04614_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10731_ (.I0(_04598_),
    .I1(\mod.u_cpu.rf_ram.memory[404][0] ),
    .S(_04614_),
    .Z(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10732_ (.I(_04615_),
    .Z(_00420_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10733_ (.I0(_04608_),
    .I1(\mod.u_cpu.rf_ram.memory[404][1] ),
    .S(_04614_),
    .Z(_04616_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10734_ (.I(_04616_),
    .Z(_00421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10735_ (.A1(_04352_),
    .A2(_04599_),
    .ZN(_04617_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10736_ (.I0(_04598_),
    .I1(\mod.u_cpu.rf_ram.memory[403][0] ),
    .S(_04617_),
    .Z(_04618_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10737_ (.I(_04618_),
    .Z(_00422_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10738_ (.I0(_04608_),
    .I1(\mod.u_cpu.rf_ram.memory[403][1] ),
    .S(_04617_),
    .Z(_04619_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10739_ (.I(_04619_),
    .Z(_00423_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10740_ (.I(_03737_),
    .Z(_04620_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10741_ (.I(_04620_),
    .Z(_04621_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10742_ (.I(_04621_),
    .Z(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10743_ (.I(_04574_),
    .Z(_04623_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10744_ (.A1(_04201_),
    .A2(_04623_),
    .ZN(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10745_ (.I0(_04622_),
    .I1(\mod.u_cpu.rf_ram.memory[402][0] ),
    .S(_04624_),
    .Z(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10746_ (.I(_04625_),
    .Z(_00424_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10747_ (.I(_04578_),
    .Z(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10748_ (.I0(_04626_),
    .I1(\mod.u_cpu.rf_ram.memory[402][1] ),
    .S(_04624_),
    .Z(_04627_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10749_ (.I(_04627_),
    .Z(_00425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10750_ (.A1(_04360_),
    .A2(_04623_),
    .ZN(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10751_ (.I0(_04622_),
    .I1(\mod.u_cpu.rf_ram.memory[401][0] ),
    .S(_04628_),
    .Z(_04629_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10752_ (.I(_04629_),
    .Z(_00426_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10753_ (.I0(_04626_),
    .I1(\mod.u_cpu.rf_ram.memory[401][1] ),
    .S(_04628_),
    .Z(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10754_ (.I(_04630_),
    .Z(_00427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10755_ (.A1(_04209_),
    .A2(_04623_),
    .ZN(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10756_ (.I0(_04622_),
    .I1(\mod.u_cpu.rf_ram.memory[400][0] ),
    .S(_04631_),
    .Z(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10757_ (.I(_04632_),
    .Z(_00428_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10758_ (.I0(_04626_),
    .I1(\mod.u_cpu.rf_ram.memory[400][1] ),
    .S(_04631_),
    .Z(_04633_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10759_ (.I(_04633_),
    .Z(_00429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10760_ (.A1(_04196_),
    .A2(_03969_),
    .ZN(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10761_ (.I0(_04622_),
    .I1(\mod.u_cpu.rf_ram.memory[3][0] ),
    .S(_04634_),
    .Z(_04635_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10762_ (.I(_04635_),
    .Z(_00430_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10763_ (.I0(_04626_),
    .I1(\mod.u_cpu.rf_ram.memory[3][1] ),
    .S(_04634_),
    .Z(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10764_ (.I(_04636_),
    .Z(_00431_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10765_ (.I(_04621_),
    .Z(_04637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10766_ (.A1(_04218_),
    .A2(_04623_),
    .ZN(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10767_ (.I0(_04637_),
    .I1(\mod.u_cpu.rf_ram.memory[398][0] ),
    .S(_04638_),
    .Z(_04639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10768_ (.I(_04639_),
    .Z(_00432_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10769_ (.I(_04496_),
    .Z(_04640_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10770_ (.I(_04640_),
    .Z(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10771_ (.I0(_04641_),
    .I1(\mod.u_cpu.rf_ram.memory[398][1] ),
    .S(_04638_),
    .Z(_04642_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10772_ (.I(_04642_),
    .Z(_00433_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10773_ (.I(_03895_),
    .Z(_04643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10774_ (.A1(_03723_),
    .A2(_04225_),
    .ZN(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10775_ (.A1(_04643_),
    .A2(_04644_),
    .ZN(_04645_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10776_ (.I0(\mod.u_cpu.rf_ram.memory[397][0] ),
    .I1(_04396_),
    .S(_04645_),
    .Z(_04646_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10777_ (.I(_04646_),
    .Z(_00434_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10778_ (.I0(\mod.u_cpu.rf_ram.memory[397][1] ),
    .I1(_04532_),
    .S(_04645_),
    .Z(_04647_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10779_ (.I(_04647_),
    .Z(_00435_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10780_ (.I(_04569_),
    .Z(_04648_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10781_ (.A1(_04233_),
    .A2(_04648_),
    .ZN(_04649_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10782_ (.I0(_04637_),
    .I1(\mod.u_cpu.rf_ram.memory[396][0] ),
    .S(_04649_),
    .Z(_04650_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10783_ (.I(_04650_),
    .Z(_00436_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10784_ (.I0(_04641_),
    .I1(\mod.u_cpu.rf_ram.memory[396][1] ),
    .S(_04649_),
    .Z(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10785_ (.I(_04651_),
    .Z(_00437_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10786_ (.A1(_04238_),
    .A2(_04648_),
    .ZN(_04652_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10787_ (.I0(_04637_),
    .I1(\mod.u_cpu.rf_ram.memory[395][0] ),
    .S(_04652_),
    .Z(_04653_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10788_ (.I(_04653_),
    .Z(_00438_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10789_ (.I0(_04641_),
    .I1(\mod.u_cpu.rf_ram.memory[395][1] ),
    .S(_04652_),
    .Z(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10790_ (.I(_04654_),
    .Z(_00439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10791_ (.A1(_04242_),
    .A2(_04648_),
    .ZN(_04655_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10792_ (.I0(_04637_),
    .I1(\mod.u_cpu.rf_ram.memory[394][0] ),
    .S(_04655_),
    .Z(_04656_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10793_ (.I(_04656_),
    .Z(_00440_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10794_ (.I0(_04641_),
    .I1(\mod.u_cpu.rf_ram.memory[394][1] ),
    .S(_04655_),
    .Z(_04657_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10795_ (.I(_04657_),
    .Z(_00441_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10796_ (.I(_03924_),
    .Z(_04658_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10797_ (.A1(_04527_),
    .A2(_04644_),
    .ZN(_04659_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10798_ (.I0(\mod.u_cpu.rf_ram.memory[393][0] ),
    .I1(_04658_),
    .S(_04659_),
    .Z(_04660_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10799_ (.I(_04660_),
    .Z(_00442_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10800_ (.I(_04531_),
    .Z(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10801_ (.I0(\mod.u_cpu.rf_ram.memory[393][1] ),
    .I1(_04661_),
    .S(_04659_),
    .Z(_04662_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10802_ (.I(_04662_),
    .Z(_00443_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10803_ (.I(_04621_),
    .Z(_04663_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10804_ (.A1(_04255_),
    .A2(_04648_),
    .ZN(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10805_ (.I0(_04663_),
    .I1(\mod.u_cpu.rf_ram.memory[392][0] ),
    .S(_04664_),
    .Z(_04665_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10806_ (.I(_04665_),
    .Z(_00444_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10807_ (.I(_04640_),
    .Z(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10808_ (.I0(_04666_),
    .I1(\mod.u_cpu.rf_ram.memory[392][1] ),
    .S(_04664_),
    .Z(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10809_ (.I(_04667_),
    .Z(_00445_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10810_ (.I(_03941_),
    .Z(_04668_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10811_ (.I(_04569_),
    .Z(_04669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10812_ (.A1(_04668_),
    .A2(_04669_),
    .ZN(_04670_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10813_ (.I0(_04663_),
    .I1(\mod.u_cpu.rf_ram.memory[391][0] ),
    .S(_04670_),
    .Z(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10814_ (.I(_04671_),
    .Z(_00446_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10815_ (.I0(_04666_),
    .I1(\mod.u_cpu.rf_ram.memory[391][1] ),
    .S(_04670_),
    .Z(_04672_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10816_ (.I(_04672_),
    .Z(_00447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10817_ (.A1(_04262_),
    .A2(_04669_),
    .ZN(_04673_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10818_ (.I0(_04663_),
    .I1(\mod.u_cpu.rf_ram.memory[390][0] ),
    .S(_04673_),
    .Z(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10819_ (.I(_04674_),
    .Z(_00448_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10820_ (.I0(_04666_),
    .I1(\mod.u_cpu.rf_ram.memory[390][1] ),
    .S(_04673_),
    .Z(_04675_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10821_ (.I(_04675_),
    .Z(_00449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10822_ (.A1(_04511_),
    .A2(_03951_),
    .ZN(_04676_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10823_ (.I0(_04663_),
    .I1(\mod.u_cpu.rf_ram.memory[38][0] ),
    .S(_04676_),
    .Z(_04677_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10824_ (.I(_04677_),
    .Z(_00450_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10825_ (.I0(_04666_),
    .I1(\mod.u_cpu.rf_ram.memory[38][1] ),
    .S(_04676_),
    .Z(_04678_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10826_ (.I(_04678_),
    .Z(_00451_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10827_ (.I(_04621_),
    .Z(_04679_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10828_ (.A1(_04272_),
    .A2(_04669_),
    .ZN(_04680_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10829_ (.I0(_04679_),
    .I1(\mod.u_cpu.rf_ram.memory[388][0] ),
    .S(_04680_),
    .Z(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10830_ (.I(_04681_),
    .Z(_00452_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10831_ (.I(_04640_),
    .Z(_04682_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10832_ (.I0(_04682_),
    .I1(\mod.u_cpu.rf_ram.memory[388][1] ),
    .S(_04680_),
    .Z(_04683_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10833_ (.I(_04683_),
    .Z(_00453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10834_ (.A1(_04277_),
    .A2(_04669_),
    .ZN(_04684_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10835_ (.I0(_04679_),
    .I1(\mod.u_cpu.rf_ram.memory[387][0] ),
    .S(_04684_),
    .Z(_04685_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10836_ (.I(_04685_),
    .Z(_00454_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10837_ (.I0(_04682_),
    .I1(\mod.u_cpu.rf_ram.memory[387][1] ),
    .S(_04684_),
    .Z(_04686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10838_ (.I(_04686_),
    .Z(_00455_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10839_ (.I(_04569_),
    .Z(_04687_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10840_ (.A1(_04281_),
    .A2(_04687_),
    .ZN(_04688_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10841_ (.I0(_04679_),
    .I1(\mod.u_cpu.rf_ram.memory[386][0] ),
    .S(_04688_),
    .Z(_04689_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10842_ (.I(_04689_),
    .Z(_00456_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10843_ (.I0(_04682_),
    .I1(\mod.u_cpu.rf_ram.memory[386][1] ),
    .S(_04688_),
    .Z(_04690_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10844_ (.I(_04690_),
    .Z(_00457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10845_ (.A1(_04285_),
    .A2(_04687_),
    .ZN(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10846_ (.I0(_04679_),
    .I1(\mod.u_cpu.rf_ram.memory[385][0] ),
    .S(_04691_),
    .Z(_04692_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10847_ (.I(_04692_),
    .Z(_00458_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10848_ (.I0(_04682_),
    .I1(\mod.u_cpu.rf_ram.memory[385][1] ),
    .S(_04691_),
    .Z(_04693_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10849_ (.I(_04693_),
    .Z(_00459_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10850_ (.I(_04620_),
    .Z(_04694_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10851_ (.I(_04694_),
    .Z(_04695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10852_ (.A1(_04290_),
    .A2(_04687_),
    .ZN(_04696_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10853_ (.I0(_04695_),
    .I1(\mod.u_cpu.rf_ram.memory[384][0] ),
    .S(_04696_),
    .Z(_04697_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10854_ (.I(_04697_),
    .Z(_00460_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10855_ (.I(_04640_),
    .Z(_04698_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10856_ (.I0(_04698_),
    .I1(\mod.u_cpu.rf_ram.memory[384][1] ),
    .S(_04696_),
    .Z(_04699_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10857_ (.I(_04699_),
    .Z(_00461_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10858_ (.I(_03990_),
    .Z(_04700_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _10859_ (.A1(\mod.u_cpu.cpu.immdec.imm11_7[3] ),
    .A2(_04222_),
    .A3(_03724_),
    .Z(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10860_ (.A1(_03992_),
    .A2(_04134_),
    .A3(_04701_),
    .ZN(_04702_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10861_ (.I(_04702_),
    .Z(_04703_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10862_ (.I(_04703_),
    .Z(_04704_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10863_ (.A1(_04700_),
    .A2(_04704_),
    .ZN(_04705_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10864_ (.A1(_04611_),
    .A2(_04705_),
    .ZN(_04706_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10865_ (.A1(_01865_),
    .A2(_04705_),
    .B(_04706_),
    .ZN(_00462_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10866_ (.I0(_04698_),
    .I1(\mod.u_cpu.rf_ram.memory[383][1] ),
    .S(_04705_),
    .Z(_04707_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10867_ (.I(_04707_),
    .Z(_00463_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10868_ (.I(_04702_),
    .Z(_04708_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10869_ (.I(_04708_),
    .Z(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10870_ (.A1(_04299_),
    .A2(_04709_),
    .ZN(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10871_ (.I0(_04695_),
    .I1(\mod.u_cpu.rf_ram.memory[382][0] ),
    .S(_04710_),
    .Z(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10872_ (.I(_04711_),
    .Z(_00464_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10873_ (.I0(_04698_),
    .I1(\mod.u_cpu.rf_ram.memory[382][1] ),
    .S(_04710_),
    .Z(_04712_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10874_ (.I(_04712_),
    .Z(_00465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10875_ (.I(_04703_),
    .Z(_04713_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10876_ (.A1(_04307_),
    .A2(_04713_),
    .ZN(_04714_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10877_ (.A1(_04611_),
    .A2(_04714_),
    .ZN(_04715_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10878_ (.A1(_01859_),
    .A2(_04714_),
    .B(_04715_),
    .ZN(_00466_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10879_ (.I0(_04698_),
    .I1(\mod.u_cpu.rf_ram.memory[381][1] ),
    .S(_04714_),
    .Z(_04716_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10880_ (.I(_04716_),
    .Z(_00467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10881_ (.A1(_04315_),
    .A2(_04709_),
    .ZN(_04717_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10882_ (.I0(_04695_),
    .I1(\mod.u_cpu.rf_ram.memory[380][0] ),
    .S(_04717_),
    .Z(_04718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10883_ (.I(_04718_),
    .Z(_00468_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10884_ (.I(_04496_),
    .Z(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10885_ (.I(_04719_),
    .Z(_04720_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10886_ (.I0(_04720_),
    .I1(\mod.u_cpu.rf_ram.memory[380][1] ),
    .S(_04717_),
    .Z(_04721_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10887_ (.I(_04721_),
    .Z(_00469_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10888_ (.A1(_04389_),
    .A2(_04108_),
    .ZN(_04722_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10889_ (.A1(_04414_),
    .A2(_04722_),
    .ZN(_04723_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10890_ (.A1(_02427_),
    .A2(_04722_),
    .B(_04723_),
    .ZN(_00470_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10891_ (.I0(\mod.u_cpu.rf_ram.memory[37][1] ),
    .I1(_04661_),
    .S(_04722_),
    .Z(_04724_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10892_ (.I(_04724_),
    .Z(_00471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10893_ (.A1(_04322_),
    .A2(_04709_),
    .ZN(_04725_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10894_ (.I0(_04695_),
    .I1(\mod.u_cpu.rf_ram.memory[378][0] ),
    .S(_04725_),
    .Z(_04726_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10895_ (.I(_04726_),
    .Z(_00472_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10896_ (.I0(_04720_),
    .I1(\mod.u_cpu.rf_ram.memory[378][1] ),
    .S(_04725_),
    .Z(_04727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10897_ (.I(_04727_),
    .Z(_00473_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10898_ (.I(_04694_),
    .Z(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10899_ (.A1(_04163_),
    .A2(_04709_),
    .ZN(_04729_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10900_ (.I0(_04728_),
    .I1(\mod.u_cpu.rf_ram.memory[377][0] ),
    .S(_04729_),
    .Z(_04730_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10901_ (.I(_04730_),
    .Z(_00474_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10902_ (.I0(_04720_),
    .I1(\mod.u_cpu.rf_ram.memory[377][1] ),
    .S(_04729_),
    .Z(_04731_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10903_ (.I(_04731_),
    .Z(_00475_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10904_ (.I(_03803_),
    .Z(_04732_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10905_ (.I(_04708_),
    .Z(_04733_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10906_ (.A1(_04732_),
    .A2(_04733_),
    .ZN(_04734_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10907_ (.I0(_04728_),
    .I1(\mod.u_cpu.rf_ram.memory[376][0] ),
    .S(_04734_),
    .Z(_04735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10908_ (.I(_04735_),
    .Z(_00476_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10909_ (.I0(_04720_),
    .I1(\mod.u_cpu.rf_ram.memory[376][1] ),
    .S(_04734_),
    .Z(_04736_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10910_ (.I(_04736_),
    .Z(_00477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10911_ (.A1(_04172_),
    .A2(_04713_),
    .ZN(_04737_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10912_ (.A1(_04611_),
    .A2(_04737_),
    .ZN(_04738_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10913_ (.A1(_01880_),
    .A2(_04737_),
    .B(_04738_),
    .ZN(_00478_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10914_ (.I(_04719_),
    .Z(_04739_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10915_ (.I0(_04739_),
    .I1(\mod.u_cpu.rf_ram.memory[375][1] ),
    .S(_04737_),
    .Z(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10916_ (.I(_04740_),
    .Z(_00479_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10917_ (.I(_03827_),
    .Z(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10918_ (.A1(_04741_),
    .A2(_04733_),
    .ZN(_04742_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10919_ (.I0(_04728_),
    .I1(\mod.u_cpu.rf_ram.memory[374][0] ),
    .S(_04742_),
    .Z(_04743_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10920_ (.I(_04743_),
    .Z(_00480_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10921_ (.I0(_04739_),
    .I1(\mod.u_cpu.rf_ram.memory[374][1] ),
    .S(_04742_),
    .Z(_04744_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10922_ (.I(_04744_),
    .Z(_00481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10923_ (.A1(_04184_),
    .A2(_04713_),
    .ZN(_04745_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10924_ (.I(_04541_),
    .Z(_04746_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10925_ (.A1(_04746_),
    .A2(_04745_),
    .ZN(_04747_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10926_ (.A1(_01876_),
    .A2(_04745_),
    .B(_04747_),
    .ZN(_00482_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10927_ (.I0(_04739_),
    .I1(\mod.u_cpu.rf_ram.memory[373][1] ),
    .S(_04745_),
    .Z(_04748_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10928_ (.I(_04748_),
    .Z(_00483_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10929_ (.I(_03841_),
    .Z(_04749_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10930_ (.A1(_04749_),
    .A2(_04733_),
    .ZN(_04750_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10931_ (.I0(_04728_),
    .I1(\mod.u_cpu.rf_ram.memory[372][0] ),
    .S(_04750_),
    .Z(_04751_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10932_ (.I(_04751_),
    .Z(_00484_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10933_ (.I0(_04739_),
    .I1(\mod.u_cpu.rf_ram.memory[372][1] ),
    .S(_04750_),
    .Z(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10934_ (.I(_04752_),
    .Z(_00485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10935_ (.I(_04694_),
    .Z(_04753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10936_ (.A1(_04352_),
    .A2(_04733_),
    .ZN(_04754_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10937_ (.I0(_04753_),
    .I1(\mod.u_cpu.rf_ram.memory[371][0] ),
    .S(_04754_),
    .Z(_04755_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10938_ (.I(_04755_),
    .Z(_00486_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10939_ (.I(_04719_),
    .Z(_04756_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10940_ (.I0(_04756_),
    .I1(\mod.u_cpu.rf_ram.memory[371][1] ),
    .S(_04754_),
    .Z(_04757_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10941_ (.I(_04757_),
    .Z(_00487_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10942_ (.I(_03857_),
    .Z(_04758_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10943_ (.I(_04708_),
    .Z(_04759_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10944_ (.A1(_04758_),
    .A2(_04759_),
    .ZN(_04760_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10945_ (.I0(_04753_),
    .I1(\mod.u_cpu.rf_ram.memory[370][0] ),
    .S(_04760_),
    .Z(_04761_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10946_ (.I(_04761_),
    .Z(_00488_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10947_ (.I0(_04756_),
    .I1(\mod.u_cpu.rf_ram.memory[370][1] ),
    .S(_04760_),
    .Z(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10948_ (.I(_04762_),
    .Z(_00489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10949_ (.A1(_04511_),
    .A2(_03961_),
    .ZN(_04763_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10950_ (.I0(_04753_),
    .I1(\mod.u_cpu.rf_ram.memory[36][0] ),
    .S(_04763_),
    .Z(_04764_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10951_ (.I(_04764_),
    .Z(_00490_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10952_ (.I0(_04756_),
    .I1(\mod.u_cpu.rf_ram.memory[36][1] ),
    .S(_04763_),
    .Z(_04765_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10953_ (.I(_04765_),
    .Z(_00491_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10954_ (.I(_03871_),
    .Z(_04766_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10955_ (.A1(_04766_),
    .A2(_04759_),
    .ZN(_04767_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10956_ (.I0(_04753_),
    .I1(\mod.u_cpu.rf_ram.memory[368][0] ),
    .S(_04767_),
    .Z(_04768_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10957_ (.I(_04768_),
    .Z(_00492_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10958_ (.I0(_04756_),
    .I1(\mod.u_cpu.rf_ram.memory[368][1] ),
    .S(_04767_),
    .Z(_04769_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10959_ (.I(_04769_),
    .Z(_00493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10960_ (.A1(_04369_),
    .A2(_04713_),
    .ZN(_04770_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10961_ (.A1(_04746_),
    .A2(_04770_),
    .ZN(_04771_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10962_ (.A1(_01897_),
    .A2(_04770_),
    .B(_04771_),
    .ZN(_00494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10963_ (.I(_04719_),
    .Z(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10964_ (.I0(_04772_),
    .I1(\mod.u_cpu.rf_ram.memory[367][1] ),
    .S(_04770_),
    .Z(_04773_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10965_ (.I(_04773_),
    .Z(_00495_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10966_ (.I(_04694_),
    .Z(_04774_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10967_ (.I(_03884_),
    .Z(_04775_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10968_ (.A1(_04775_),
    .A2(_04759_),
    .ZN(_04776_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10969_ (.I0(_04774_),
    .I1(\mod.u_cpu.rf_ram.memory[366][0] ),
    .S(_04776_),
    .Z(_04777_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10970_ (.I(_04777_),
    .Z(_00496_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10971_ (.I0(_04772_),
    .I1(\mod.u_cpu.rf_ram.memory[366][1] ),
    .S(_04776_),
    .Z(_04778_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10972_ (.I(_04778_),
    .Z(_00497_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _10973_ (.A1(_03663_),
    .A2(_04223_),
    .A3(_03724_),
    .ZN(_04779_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10974_ (.A1(_04227_),
    .A2(_04779_),
    .ZN(_04780_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10975_ (.A1(_04377_),
    .A2(_04780_),
    .ZN(_04781_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10976_ (.A1(_04414_),
    .A2(_04781_),
    .ZN(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10977_ (.A1(_01894_),
    .A2(_04781_),
    .B(_04782_),
    .ZN(_00498_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10978_ (.I0(\mod.u_cpu.rf_ram.memory[365][1] ),
    .I1(_04661_),
    .S(_04781_),
    .Z(_04783_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10979_ (.I(_04783_),
    .Z(_00499_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10980_ (.I(_03903_),
    .Z(_04784_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10981_ (.A1(_04784_),
    .A2(_04759_),
    .ZN(_04785_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10982_ (.I0(_04774_),
    .I1(\mod.u_cpu.rf_ram.memory[364][0] ),
    .S(_04785_),
    .Z(_04786_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10983_ (.I(_04786_),
    .Z(_00500_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10984_ (.I0(_04772_),
    .I1(\mod.u_cpu.rf_ram.memory[364][1] ),
    .S(_04785_),
    .Z(_04787_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10985_ (.I(_04787_),
    .Z(_00501_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10986_ (.I(_04703_),
    .Z(_04788_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10987_ (.A1(_04238_),
    .A2(_04788_),
    .ZN(_04789_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10988_ (.I0(_04774_),
    .I1(\mod.u_cpu.rf_ram.memory[363][0] ),
    .S(_04789_),
    .Z(_04790_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10989_ (.I(_04790_),
    .Z(_00502_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10990_ (.I0(_04772_),
    .I1(\mod.u_cpu.rf_ram.memory[363][1] ),
    .S(_04789_),
    .Z(_04791_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10991_ (.I(_04791_),
    .Z(_00503_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10992_ (.I(_03917_),
    .Z(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10993_ (.A1(_04792_),
    .A2(_04788_),
    .ZN(_04793_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10994_ (.I0(_04774_),
    .I1(\mod.u_cpu.rf_ram.memory[362][0] ),
    .S(_04793_),
    .Z(_04794_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10995_ (.I(_04794_),
    .Z(_00504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10996_ (.I(_03761_),
    .Z(_04795_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10997_ (.I(_04795_),
    .Z(_04796_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10998_ (.I(_04796_),
    .Z(_04797_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10999_ (.I0(_04797_),
    .I1(\mod.u_cpu.rf_ram.memory[362][1] ),
    .S(_04793_),
    .Z(_04798_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11000_ (.I(_04798_),
    .Z(_00505_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11001_ (.A1(_04527_),
    .A2(_04780_),
    .ZN(_04799_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11002_ (.I0(\mod.u_cpu.rf_ram.memory[361][0] ),
    .I1(_04658_),
    .S(_04799_),
    .Z(_04800_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11003_ (.I(_04800_),
    .Z(_00506_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11004_ (.I0(\mod.u_cpu.rf_ram.memory[361][1] ),
    .I1(_04661_),
    .S(_04799_),
    .Z(_04801_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11005_ (.I(_04801_),
    .Z(_00507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11006_ (.I(_04620_),
    .Z(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11007_ (.I(_04802_),
    .Z(_04803_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11008_ (.I(_03931_),
    .Z(_04804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11009_ (.A1(_04804_),
    .A2(_04788_),
    .ZN(_04805_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11010_ (.I0(_04803_),
    .I1(\mod.u_cpu.rf_ram.memory[360][0] ),
    .S(_04805_),
    .Z(_04806_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11011_ (.I(_04806_),
    .Z(_00508_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11012_ (.I0(_04797_),
    .I1(\mod.u_cpu.rf_ram.memory[360][1] ),
    .S(_04805_),
    .Z(_04807_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11013_ (.I(_04807_),
    .Z(_00509_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11014_ (.I(_04250_),
    .Z(_04808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11015_ (.A1(_04808_),
    .A2(_03969_),
    .ZN(_04809_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11016_ (.I0(_04803_),
    .I1(\mod.u_cpu.rf_ram.memory[35][0] ),
    .S(_04809_),
    .Z(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11017_ (.I(_04810_),
    .Z(_00510_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11018_ (.I0(_04797_),
    .I1(\mod.u_cpu.rf_ram.memory[35][1] ),
    .S(_04809_),
    .Z(_04811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11019_ (.I(_04811_),
    .Z(_00511_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11020_ (.I(_03949_),
    .Z(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11021_ (.A1(_04812_),
    .A2(_04788_),
    .ZN(_04813_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11022_ (.I0(_04803_),
    .I1(\mod.u_cpu.rf_ram.memory[358][0] ),
    .S(_04813_),
    .Z(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11023_ (.I(_04814_),
    .Z(_00512_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11024_ (.I0(_04797_),
    .I1(\mod.u_cpu.rf_ram.memory[358][1] ),
    .S(_04813_),
    .Z(_04815_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11025_ (.I(_04815_),
    .Z(_00513_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11026_ (.A1(_04412_),
    .A2(_04780_),
    .ZN(_04816_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11027_ (.I(_03898_),
    .Z(_04817_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11028_ (.A1(_04817_),
    .A2(_04816_),
    .ZN(_04818_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11029_ (.A1(_01903_),
    .A2(_04816_),
    .B(_04818_),
    .ZN(_00514_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11030_ (.I(_04531_),
    .Z(_04819_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11031_ (.I0(\mod.u_cpu.rf_ram.memory[357][1] ),
    .I1(_04819_),
    .S(_04816_),
    .Z(_04820_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11032_ (.I(_04820_),
    .Z(_00515_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11033_ (.I(_03959_),
    .Z(_04821_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11034_ (.I(_04703_),
    .Z(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11035_ (.A1(_04821_),
    .A2(_04822_),
    .ZN(_04823_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11036_ (.I0(_04803_),
    .I1(\mod.u_cpu.rf_ram.memory[356][0] ),
    .S(_04823_),
    .Z(_04824_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11037_ (.I(_04824_),
    .Z(_00516_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11038_ (.I(_04796_),
    .Z(_04825_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11039_ (.I0(_04825_),
    .I1(\mod.u_cpu.rf_ram.memory[356][1] ),
    .S(_04823_),
    .Z(_04826_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11040_ (.I(_04826_),
    .Z(_00517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11041_ (.I(_04802_),
    .Z(_04827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11042_ (.A1(_04277_),
    .A2(_04822_),
    .ZN(_04828_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11043_ (.I0(_04827_),
    .I1(\mod.u_cpu.rf_ram.memory[355][0] ),
    .S(_04828_),
    .Z(_04829_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11044_ (.I(_04829_),
    .Z(_00518_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11045_ (.I0(_04825_),
    .I1(\mod.u_cpu.rf_ram.memory[355][1] ),
    .S(_04828_),
    .Z(_04830_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11046_ (.I(_04830_),
    .Z(_00519_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11047_ (.I(_03973_),
    .Z(_04831_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11048_ (.A1(_04831_),
    .A2(_04822_),
    .ZN(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11049_ (.I0(_04827_),
    .I1(\mod.u_cpu.rf_ram.memory[354][0] ),
    .S(_04832_),
    .Z(_04833_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11050_ (.I(_04833_),
    .Z(_00520_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11051_ (.I0(_04825_),
    .I1(\mod.u_cpu.rf_ram.memory[354][1] ),
    .S(_04832_),
    .Z(_04834_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11052_ (.I(_04834_),
    .Z(_00521_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11053_ (.A1(_04285_),
    .A2(_04822_),
    .ZN(_04835_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11054_ (.I0(_04827_),
    .I1(\mod.u_cpu.rf_ram.memory[353][0] ),
    .S(_04835_),
    .Z(_04836_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11055_ (.I(_04836_),
    .Z(_00522_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11056_ (.I0(_04825_),
    .I1(\mod.u_cpu.rf_ram.memory[353][1] ),
    .S(_04835_),
    .Z(_04837_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11057_ (.I(_04837_),
    .Z(_00523_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11058_ (.I(_03984_),
    .Z(_04838_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11059_ (.A1(_04838_),
    .A2(_04704_),
    .ZN(_04839_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11060_ (.I0(_04827_),
    .I1(\mod.u_cpu.rf_ram.memory[352][0] ),
    .S(_04839_),
    .Z(_04840_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11061_ (.I(_04840_),
    .Z(_00524_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11062_ (.I(_04796_),
    .Z(_04841_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11063_ (.I0(_04841_),
    .I1(\mod.u_cpu.rf_ram.memory[352][1] ),
    .S(_04839_),
    .Z(_04842_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11064_ (.I(_04842_),
    .Z(_00525_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11065_ (.I(_04802_),
    .Z(_04843_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11066_ (.I(_03990_),
    .Z(_04844_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11067_ (.I(_04844_),
    .Z(_04845_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11068_ (.A1(_04300_),
    .A2(_04701_),
    .ZN(_04846_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11069_ (.I(_04846_),
    .Z(_04847_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11070_ (.I(_04847_),
    .Z(_04848_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11071_ (.A1(_04845_),
    .A2(_04848_),
    .ZN(_04849_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11072_ (.I0(_04843_),
    .I1(\mod.u_cpu.rf_ram.memory[351][0] ),
    .S(_04849_),
    .Z(_04850_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11073_ (.I(_04850_),
    .Z(_00526_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11074_ (.I0(_04841_),
    .I1(\mod.u_cpu.rf_ram.memory[351][1] ),
    .S(_04849_),
    .Z(_04851_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11075_ (.I(_04851_),
    .Z(_00527_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11076_ (.I(_03750_),
    .Z(_04852_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11077_ (.A1(_04852_),
    .A2(_04848_),
    .ZN(_04853_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11078_ (.I0(_04843_),
    .I1(\mod.u_cpu.rf_ram.memory[350][0] ),
    .S(_04853_),
    .Z(_04854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11079_ (.I(_04854_),
    .Z(_00528_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11080_ (.I0(_04841_),
    .I1(\mod.u_cpu.rf_ram.memory[350][1] ),
    .S(_04853_),
    .Z(_04855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11081_ (.I(_04855_),
    .Z(_00529_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11082_ (.A1(_04808_),
    .A2(_03975_),
    .ZN(_04856_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11083_ (.I0(_04843_),
    .I1(\mod.u_cpu.rf_ram.memory[34][0] ),
    .S(_04856_),
    .Z(_04857_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11084_ (.I(_04857_),
    .Z(_00530_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11085_ (.I0(_04841_),
    .I1(\mod.u_cpu.rf_ram.memory[34][1] ),
    .S(_04856_),
    .Z(_04858_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11086_ (.I(_04858_),
    .Z(_00531_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11087_ (.I(_03780_),
    .Z(_04859_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11088_ (.A1(_04859_),
    .A2(_04848_),
    .ZN(_04860_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11089_ (.I0(_04843_),
    .I1(\mod.u_cpu.rf_ram.memory[348][0] ),
    .S(_04860_),
    .Z(_04861_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11090_ (.I(_04861_),
    .Z(_00532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11091_ (.I(_04796_),
    .Z(_04862_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11092_ (.I0(_04862_),
    .I1(\mod.u_cpu.rf_ram.memory[348][1] ),
    .S(_04860_),
    .Z(_04863_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11093_ (.I(_04863_),
    .Z(_00533_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11094_ (.I(_04802_),
    .Z(_04864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11095_ (.A1(_04457_),
    .A2(_04848_),
    .ZN(_04865_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11096_ (.I0(_04864_),
    .I1(\mod.u_cpu.rf_ram.memory[347][0] ),
    .S(_04865_),
    .Z(_04866_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11097_ (.I(_04866_),
    .Z(_00534_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11098_ (.I0(_04862_),
    .I1(\mod.u_cpu.rf_ram.memory[347][1] ),
    .S(_04865_),
    .Z(_04867_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11099_ (.I(_04867_),
    .Z(_00535_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11100_ (.I(_03795_),
    .Z(_04868_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11101_ (.I(_04847_),
    .Z(_04869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11102_ (.A1(_04868_),
    .A2(_04869_),
    .ZN(_04870_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11103_ (.I0(_04864_),
    .I1(\mod.u_cpu.rf_ram.memory[346][0] ),
    .S(_04870_),
    .Z(_04871_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11104_ (.I(_04871_),
    .Z(_00536_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11105_ (.I0(_04862_),
    .I1(\mod.u_cpu.rf_ram.memory[346][1] ),
    .S(_04870_),
    .Z(_04872_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11106_ (.I(_04872_),
    .Z(_00537_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11107_ (.I(_04024_),
    .Z(_04873_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11108_ (.A1(_04873_),
    .A2(_04869_),
    .ZN(_04874_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11109_ (.I0(_04864_),
    .I1(\mod.u_cpu.rf_ram.memory[345][0] ),
    .S(_04874_),
    .Z(_04875_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11110_ (.I(_04875_),
    .Z(_00538_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11111_ (.I0(_04862_),
    .I1(\mod.u_cpu.rf_ram.memory[345][1] ),
    .S(_04874_),
    .Z(_04876_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11112_ (.I(_04876_),
    .Z(_00539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11113_ (.A1(_04732_),
    .A2(_04869_),
    .ZN(_04877_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11114_ (.I0(_04864_),
    .I1(\mod.u_cpu.rf_ram.memory[344][0] ),
    .S(_04877_),
    .Z(_04878_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11115_ (.I(_04878_),
    .Z(_00540_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11116_ (.I(_04795_),
    .Z(_04879_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11117_ (.I(_04879_),
    .Z(_04880_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11118_ (.I0(_04880_),
    .I1(\mod.u_cpu.rf_ram.memory[344][1] ),
    .S(_04877_),
    .Z(_04881_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11119_ (.I(_04881_),
    .Z(_00541_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11120_ (.I(_04620_),
    .Z(_04882_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11121_ (.I(_04882_),
    .Z(_04883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11122_ (.A1(_03879_),
    .A2(_04869_),
    .ZN(_04884_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11123_ (.I0(_04883_),
    .I1(\mod.u_cpu.rf_ram.memory[343][0] ),
    .S(_04884_),
    .Z(_04885_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11124_ (.I(_04885_),
    .Z(_00542_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11125_ (.I0(_04880_),
    .I1(\mod.u_cpu.rf_ram.memory[343][1] ),
    .S(_04884_),
    .Z(_04886_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11126_ (.I(_04886_),
    .Z(_00543_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11127_ (.I(_04847_),
    .Z(_04887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11128_ (.A1(_04741_),
    .A2(_04887_),
    .ZN(_04888_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11129_ (.I0(_04883_),
    .I1(\mod.u_cpu.rf_ram.memory[342][0] ),
    .S(_04888_),
    .Z(_04889_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11130_ (.I(_04889_),
    .Z(_00544_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11131_ (.I0(_04880_),
    .I1(\mod.u_cpu.rf_ram.memory[342][1] ),
    .S(_04888_),
    .Z(_04890_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11132_ (.I(_04890_),
    .Z(_00545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11133_ (.A1(_04014_),
    .A2(_04887_),
    .ZN(_04891_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11134_ (.I0(_04883_),
    .I1(\mod.u_cpu.rf_ram.memory[341][0] ),
    .S(_04891_),
    .Z(_04892_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11135_ (.I(_04892_),
    .Z(_00546_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11136_ (.I0(_04880_),
    .I1(\mod.u_cpu.rf_ram.memory[341][1] ),
    .S(_04891_),
    .Z(_04893_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11137_ (.I(_04893_),
    .Z(_00547_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11138_ (.A1(_04749_),
    .A2(_04887_),
    .ZN(_04894_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11139_ (.I0(_04883_),
    .I1(\mod.u_cpu.rf_ram.memory[340][0] ),
    .S(_04894_),
    .Z(_04895_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11140_ (.I(_04895_),
    .Z(_00548_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11141_ (.I(_04879_),
    .Z(_04896_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11142_ (.I0(_04896_),
    .I1(\mod.u_cpu.rf_ram.memory[340][1] ),
    .S(_04894_),
    .Z(_04897_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11143_ (.I(_04897_),
    .Z(_00549_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11144_ (.A1(_03809_),
    .A2(_03980_),
    .Z(_04898_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11145_ (.I0(\mod.u_cpu.rf_ram.memory[33][0] ),
    .I1(_04658_),
    .S(_04898_),
    .Z(_04899_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11146_ (.I(_04899_),
    .Z(_00550_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11147_ (.I0(\mod.u_cpu.rf_ram.memory[33][1] ),
    .I1(_04819_),
    .S(_04898_),
    .Z(_04900_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11148_ (.I(_04900_),
    .Z(_00551_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11149_ (.I(_04882_),
    .Z(_04901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11150_ (.A1(_04758_),
    .A2(_04887_),
    .ZN(_04902_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11151_ (.I0(_04901_),
    .I1(\mod.u_cpu.rf_ram.memory[338][0] ),
    .S(_04902_),
    .Z(_04903_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11152_ (.I(_04903_),
    .Z(_00552_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11153_ (.I0(_04896_),
    .I1(\mod.u_cpu.rf_ram.memory[338][1] ),
    .S(_04902_),
    .Z(_04904_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11154_ (.I(_04904_),
    .Z(_00553_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11155_ (.I(_04846_),
    .Z(_04905_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11156_ (.I(_04905_),
    .Z(_04906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11157_ (.A1(_04360_),
    .A2(_04906_),
    .ZN(_04907_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11158_ (.I0(_04901_),
    .I1(\mod.u_cpu.rf_ram.memory[337][0] ),
    .S(_04907_),
    .Z(_04908_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11159_ (.I(_04908_),
    .Z(_00554_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11160_ (.I0(_04896_),
    .I1(\mod.u_cpu.rf_ram.memory[337][1] ),
    .S(_04907_),
    .Z(_04909_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11161_ (.I(_04909_),
    .Z(_00555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11162_ (.A1(_04766_),
    .A2(_04906_),
    .ZN(_04910_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11163_ (.I0(_04901_),
    .I1(\mod.u_cpu.rf_ram.memory[336][0] ),
    .S(_04910_),
    .Z(_04911_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11164_ (.I(_04911_),
    .Z(_00556_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11165_ (.I0(_04896_),
    .I1(\mod.u_cpu.rf_ram.memory[336][1] ),
    .S(_04910_),
    .Z(_04912_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11166_ (.I(_04912_),
    .Z(_00557_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11167_ (.I(_04067_),
    .Z(_04913_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11168_ (.A1(_04913_),
    .A2(_04906_),
    .ZN(_04914_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11169_ (.I0(_04901_),
    .I1(\mod.u_cpu.rf_ram.memory[335][0] ),
    .S(_04914_),
    .Z(_04915_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11170_ (.I(_04915_),
    .Z(_00558_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11171_ (.I(_04879_),
    .Z(_04916_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11172_ (.I0(_04916_),
    .I1(\mod.u_cpu.rf_ram.memory[335][1] ),
    .S(_04914_),
    .Z(_04917_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11173_ (.I(_04917_),
    .Z(_00559_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11174_ (.I(_04882_),
    .Z(_04918_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11175_ (.A1(_04775_),
    .A2(_04906_),
    .ZN(_04919_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11176_ (.I0(_04918_),
    .I1(\mod.u_cpu.rf_ram.memory[334][0] ),
    .S(_04919_),
    .Z(_04920_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11177_ (.I(_04920_),
    .Z(_00560_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11178_ (.I0(_04916_),
    .I1(\mod.u_cpu.rf_ram.memory[334][1] ),
    .S(_04919_),
    .Z(_04921_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11179_ (.I(_04921_),
    .Z(_00561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11180_ (.A1(_04379_),
    .A2(_04779_),
    .ZN(_04922_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11181_ (.A1(_04643_),
    .A2(_04922_),
    .ZN(_04923_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11182_ (.I0(\mod.u_cpu.rf_ram.memory[333][0] ),
    .I1(_04658_),
    .S(_04923_),
    .Z(_04924_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11183_ (.I(_04924_),
    .Z(_00562_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11184_ (.I0(\mod.u_cpu.rf_ram.memory[333][1] ),
    .I1(_04819_),
    .S(_04923_),
    .Z(_04925_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11185_ (.I(_04925_),
    .Z(_00563_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11186_ (.I(_04905_),
    .Z(_04926_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11187_ (.A1(_04784_),
    .A2(_04926_),
    .ZN(_04927_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11188_ (.I0(_04918_),
    .I1(\mod.u_cpu.rf_ram.memory[332][0] ),
    .S(_04927_),
    .Z(_04928_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11189_ (.I(_04928_),
    .Z(_00564_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11190_ (.I0(_04916_),
    .I1(\mod.u_cpu.rf_ram.memory[332][1] ),
    .S(_04927_),
    .Z(_04929_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11191_ (.I(_04929_),
    .Z(_00565_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11192_ (.I(_03909_),
    .Z(_04930_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11193_ (.A1(_04930_),
    .A2(_04926_),
    .ZN(_04931_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11194_ (.I0(_04918_),
    .I1(\mod.u_cpu.rf_ram.memory[331][0] ),
    .S(_04931_),
    .Z(_04932_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11195_ (.I(_04932_),
    .Z(_00566_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11196_ (.I0(_04916_),
    .I1(\mod.u_cpu.rf_ram.memory[331][1] ),
    .S(_04931_),
    .Z(_04933_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11197_ (.I(_04933_),
    .Z(_00567_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11198_ (.A1(_04792_),
    .A2(_04926_),
    .ZN(_04934_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11199_ (.I0(_04918_),
    .I1(\mod.u_cpu.rf_ram.memory[330][0] ),
    .S(_04934_),
    .Z(_04935_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11200_ (.I(_04935_),
    .Z(_00568_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11201_ (.I(_04879_),
    .Z(_04936_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11202_ (.I0(_04936_),
    .I1(\mod.u_cpu.rf_ram.memory[330][1] ),
    .S(_04934_),
    .Z(_04937_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11203_ (.I(_04937_),
    .Z(_00569_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11204_ (.I(_04882_),
    .Z(_04938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11205_ (.A1(_04808_),
    .A2(_03986_),
    .ZN(_04939_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11206_ (.I0(_04938_),
    .I1(\mod.u_cpu.rf_ram.memory[32][0] ),
    .S(_04939_),
    .Z(_04940_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11207_ (.I(_04940_),
    .Z(_00570_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11208_ (.I0(_04936_),
    .I1(\mod.u_cpu.rf_ram.memory[32][1] ),
    .S(_04939_),
    .Z(_04941_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11209_ (.I(_04941_),
    .Z(_00571_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11210_ (.A1(_04804_),
    .A2(_04926_),
    .ZN(_04942_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11211_ (.I0(_04938_),
    .I1(\mod.u_cpu.rf_ram.memory[328][0] ),
    .S(_04942_),
    .Z(_04943_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11212_ (.I(_04943_),
    .Z(_00572_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11213_ (.I0(_04936_),
    .I1(\mod.u_cpu.rf_ram.memory[328][1] ),
    .S(_04942_),
    .Z(_04944_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11214_ (.I(_04944_),
    .Z(_00573_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11215_ (.I(_04905_),
    .Z(_04945_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11216_ (.A1(_04668_),
    .A2(_04945_),
    .ZN(_04946_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11217_ (.I0(_04938_),
    .I1(\mod.u_cpu.rf_ram.memory[327][0] ),
    .S(_04946_),
    .Z(_04947_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11218_ (.I(_04947_),
    .Z(_00574_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11219_ (.I0(_04936_),
    .I1(\mod.u_cpu.rf_ram.memory[327][1] ),
    .S(_04946_),
    .Z(_04948_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11220_ (.I(_04948_),
    .Z(_00575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11221_ (.A1(_04812_),
    .A2(_04945_),
    .ZN(_04949_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11222_ (.I0(_04938_),
    .I1(\mod.u_cpu.rf_ram.memory[326][0] ),
    .S(_04949_),
    .Z(_04950_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11223_ (.I(_04950_),
    .Z(_00576_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11224_ (.I(_04795_),
    .Z(_04951_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11225_ (.I(_04951_),
    .Z(_04952_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11226_ (.I0(_04952_),
    .I1(\mod.u_cpu.rf_ram.memory[326][1] ),
    .S(_04949_),
    .Z(_04953_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11227_ (.I(_04953_),
    .Z(_00577_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11228_ (.I(_03924_),
    .Z(_04954_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11229_ (.I(_04107_),
    .Z(_04955_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11230_ (.A1(_04955_),
    .A2(_04922_),
    .ZN(_04956_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11231_ (.I0(\mod.u_cpu.rf_ram.memory[325][0] ),
    .I1(_04954_),
    .S(_04956_),
    .Z(_04957_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11232_ (.I(_04957_),
    .Z(_00578_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11233_ (.I0(\mod.u_cpu.rf_ram.memory[325][1] ),
    .I1(_04819_),
    .S(_04956_),
    .Z(_04958_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11234_ (.I(_04958_),
    .Z(_00579_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11235_ (.I(_03737_),
    .Z(_04959_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11236_ (.I(_04959_),
    .Z(_04960_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11237_ (.I(_04960_),
    .Z(_04961_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11238_ (.A1(_04821_),
    .A2(_04945_),
    .ZN(_04962_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11239_ (.I0(_04961_),
    .I1(\mod.u_cpu.rf_ram.memory[324][0] ),
    .S(_04962_),
    .Z(_04963_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11240_ (.I(_04963_),
    .Z(_00580_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11241_ (.I0(_04952_),
    .I1(\mod.u_cpu.rf_ram.memory[324][1] ),
    .S(_04962_),
    .Z(_04964_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11242_ (.I(_04964_),
    .Z(_00581_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11243_ (.I(_03967_),
    .Z(_04965_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11244_ (.A1(_04965_),
    .A2(_04945_),
    .ZN(_04966_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11245_ (.I0(_04961_),
    .I1(\mod.u_cpu.rf_ram.memory[323][0] ),
    .S(_04966_),
    .Z(_04967_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11246_ (.I(_04967_),
    .Z(_00582_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11247_ (.I0(_04952_),
    .I1(\mod.u_cpu.rf_ram.memory[323][1] ),
    .S(_04966_),
    .Z(_04968_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11248_ (.I(_04968_),
    .Z(_00583_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11249_ (.I(_04905_),
    .Z(_04969_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11250_ (.A1(_04831_),
    .A2(_04969_),
    .ZN(_04970_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11251_ (.I0(_04961_),
    .I1(\mod.u_cpu.rf_ram.memory[322][0] ),
    .S(_04970_),
    .Z(_04971_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11252_ (.I(_04971_),
    .Z(_00584_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11253_ (.I0(_04952_),
    .I1(\mod.u_cpu.rf_ram.memory[322][1] ),
    .S(_04970_),
    .Z(_04972_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11254_ (.I(_04972_),
    .Z(_00585_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11255_ (.I(_04125_),
    .Z(_04973_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11256_ (.A1(_04973_),
    .A2(_04969_),
    .ZN(_04974_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11257_ (.I0(_04961_),
    .I1(\mod.u_cpu.rf_ram.memory[321][0] ),
    .S(_04974_),
    .Z(_04975_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11258_ (.I(_04975_),
    .Z(_00586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11259_ (.I(_04951_),
    .Z(_04976_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11260_ (.I0(_04976_),
    .I1(\mod.u_cpu.rf_ram.memory[321][1] ),
    .S(_04974_),
    .Z(_04977_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11261_ (.I(_04977_),
    .Z(_00587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11262_ (.I(_04960_),
    .Z(_04978_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11263_ (.A1(_04838_),
    .A2(_04969_),
    .ZN(_04979_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11264_ (.I0(_04978_),
    .I1(\mod.u_cpu.rf_ram.memory[320][0] ),
    .S(_04979_),
    .Z(_04980_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11265_ (.I(_04980_),
    .Z(_00588_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11266_ (.I0(_04976_),
    .I1(\mod.u_cpu.rf_ram.memory[320][1] ),
    .S(_04979_),
    .Z(_04981_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11267_ (.I(_04981_),
    .Z(_00589_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11268_ (.I(_04194_),
    .Z(_04982_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11269_ (.I(_04982_),
    .Z(_04983_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11270_ (.I(_04844_),
    .Z(_04984_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11271_ (.A1(_04983_),
    .A2(_04984_),
    .ZN(_04985_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11272_ (.A1(_04746_),
    .A2(_04985_),
    .ZN(_04986_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11273_ (.A1(_02398_),
    .A2(_04985_),
    .B(_04986_),
    .ZN(_00590_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11274_ (.I0(_04976_),
    .I1(\mod.u_cpu.rf_ram.memory[31][1] ),
    .S(_04985_),
    .Z(_04987_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11275_ (.I(_04987_),
    .Z(_00591_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11276_ (.A1(_03755_),
    .A2(_04701_),
    .ZN(_04988_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11277_ (.I(_04988_),
    .Z(_04989_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11278_ (.I(_04989_),
    .Z(_04990_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11279_ (.A1(_04852_),
    .A2(_04990_),
    .ZN(_04991_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11280_ (.I0(_04978_),
    .I1(\mod.u_cpu.rf_ram.memory[318][0] ),
    .S(_04991_),
    .Z(_04992_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11281_ (.I(_04992_),
    .Z(_00592_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11282_ (.I0(_04976_),
    .I1(\mod.u_cpu.rf_ram.memory[318][1] ),
    .S(_04991_),
    .Z(_04993_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11283_ (.I(_04993_),
    .Z(_00593_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11284_ (.I(_03769_),
    .Z(_04994_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11285_ (.I(_04988_),
    .Z(_04995_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11286_ (.I(_04995_),
    .Z(_04996_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11287_ (.A1(_04994_),
    .A2(_04996_),
    .ZN(_04997_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11288_ (.A1(_04746_),
    .A2(_04997_),
    .ZN(_04998_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11289_ (.A1(_01921_),
    .A2(_04997_),
    .B(_04998_),
    .ZN(_00594_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11290_ (.I(_04951_),
    .Z(_04999_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11291_ (.I0(_04999_),
    .I1(\mod.u_cpu.rf_ram.memory[317][1] ),
    .S(_04997_),
    .Z(_05000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11292_ (.I(_05000_),
    .Z(_00595_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11293_ (.A1(_04859_),
    .A2(_04990_),
    .ZN(_05001_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11294_ (.I0(_04978_),
    .I1(\mod.u_cpu.rf_ram.memory[316][0] ),
    .S(_05001_),
    .Z(_05002_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11295_ (.I(_05002_),
    .Z(_00596_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11296_ (.I0(_04999_),
    .I1(\mod.u_cpu.rf_ram.memory[316][1] ),
    .S(_05001_),
    .Z(_05003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11297_ (.I(_05003_),
    .Z(_00597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11298_ (.A1(_04457_),
    .A2(_04990_),
    .ZN(_05004_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11299_ (.I0(_04978_),
    .I1(\mod.u_cpu.rf_ram.memory[315][0] ),
    .S(_05004_),
    .Z(_05005_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11300_ (.I(_05005_),
    .Z(_00598_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11301_ (.I0(_04999_),
    .I1(\mod.u_cpu.rf_ram.memory[315][1] ),
    .S(_05004_),
    .Z(_05006_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11302_ (.I(_05006_),
    .Z(_00599_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11303_ (.I(_04960_),
    .Z(_05007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11304_ (.A1(_04868_),
    .A2(_04990_),
    .ZN(_05008_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11305_ (.I0(_05007_),
    .I1(\mod.u_cpu.rf_ram.memory[314][0] ),
    .S(_05008_),
    .Z(_05009_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11306_ (.I(_05009_),
    .Z(_00600_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11307_ (.I0(_04999_),
    .I1(\mod.u_cpu.rf_ram.memory[314][1] ),
    .S(_05008_),
    .Z(_05010_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11308_ (.I(_05010_),
    .Z(_00601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11309_ (.I(_04989_),
    .Z(_05011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11310_ (.A1(_04873_),
    .A2(_05011_),
    .ZN(_05012_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11311_ (.I0(_05007_),
    .I1(\mod.u_cpu.rf_ram.memory[313][0] ),
    .S(_05012_),
    .Z(_05013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11312_ (.I(_05013_),
    .Z(_00602_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11313_ (.I(_04951_),
    .Z(_05014_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11314_ (.I0(_05014_),
    .I1(\mod.u_cpu.rf_ram.memory[313][1] ),
    .S(_05012_),
    .Z(_05015_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11315_ (.I(_05015_),
    .Z(_00603_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11316_ (.A1(_04732_),
    .A2(_05011_),
    .ZN(_05016_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11317_ (.I0(_05007_),
    .I1(\mod.u_cpu.rf_ram.memory[312][0] ),
    .S(_05016_),
    .Z(_05017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11318_ (.I(_05017_),
    .Z(_00604_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11319_ (.I0(_05014_),
    .I1(\mod.u_cpu.rf_ram.memory[312][1] ),
    .S(_05016_),
    .Z(_05018_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11320_ (.I(_05018_),
    .Z(_00605_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11321_ (.I(_03821_),
    .Z(_05019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11322_ (.I(_04995_),
    .Z(_05020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11323_ (.A1(_05019_),
    .A2(_05020_),
    .ZN(_05021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11324_ (.I(_04541_),
    .Z(_05022_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11325_ (.A1(_05022_),
    .A2(_05021_),
    .ZN(_05023_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11326_ (.A1(_01939_),
    .A2(_05021_),
    .B(_05023_),
    .ZN(_00606_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11327_ (.I0(_05014_),
    .I1(\mod.u_cpu.rf_ram.memory[311][1] ),
    .S(_05021_),
    .Z(_05024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11328_ (.I(_05024_),
    .Z(_00607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11329_ (.A1(_04741_),
    .A2(_05011_),
    .ZN(_05025_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11330_ (.I0(_05007_),
    .I1(\mod.u_cpu.rf_ram.memory[310][0] ),
    .S(_05025_),
    .Z(_05026_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11331_ (.I(_05026_),
    .Z(_00608_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11332_ (.I0(_05014_),
    .I1(\mod.u_cpu.rf_ram.memory[310][1] ),
    .S(_05025_),
    .Z(_05027_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11333_ (.I(_05027_),
    .Z(_00609_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11334_ (.I(_04960_),
    .Z(_05028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11335_ (.A1(_04196_),
    .A2(_03752_),
    .ZN(_05029_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11336_ (.I0(_05028_),
    .I1(\mod.u_cpu.rf_ram.memory[30][0] ),
    .S(_05029_),
    .Z(_05030_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11337_ (.I(_05030_),
    .Z(_00610_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11338_ (.I(_04795_),
    .Z(_05031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11339_ (.I(_05031_),
    .Z(_05032_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11340_ (.I0(_05032_),
    .I1(\mod.u_cpu.rf_ram.memory[30][1] ),
    .S(_05029_),
    .Z(_05033_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11341_ (.I(_05033_),
    .Z(_00611_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11342_ (.A1(_04749_),
    .A2(_05011_),
    .ZN(_05034_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11343_ (.I0(_05028_),
    .I1(\mod.u_cpu.rf_ram.memory[308][0] ),
    .S(_05034_),
    .Z(_05035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11344_ (.I(_05035_),
    .Z(_00612_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11345_ (.I0(_05032_),
    .I1(\mod.u_cpu.rf_ram.memory[308][1] ),
    .S(_05034_),
    .Z(_05036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11346_ (.I(_05036_),
    .Z(_00613_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11347_ (.I(_03849_),
    .Z(_05037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11348_ (.I(_04989_),
    .Z(_05038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11349_ (.A1(_05037_),
    .A2(_05038_),
    .ZN(_05039_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11350_ (.I0(_05028_),
    .I1(\mod.u_cpu.rf_ram.memory[307][0] ),
    .S(_05039_),
    .Z(_05040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11351_ (.I(_05040_),
    .Z(_00614_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11352_ (.I0(_05032_),
    .I1(\mod.u_cpu.rf_ram.memory[307][1] ),
    .S(_05039_),
    .Z(_05041_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11353_ (.I(_05041_),
    .Z(_00615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11354_ (.A1(_04758_),
    .A2(_05038_),
    .ZN(_05042_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11355_ (.I0(_05028_),
    .I1(\mod.u_cpu.rf_ram.memory[306][0] ),
    .S(_05042_),
    .Z(_05043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11356_ (.I(_05043_),
    .Z(_00616_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11357_ (.I0(_05032_),
    .I1(\mod.u_cpu.rf_ram.memory[306][1] ),
    .S(_05042_),
    .Z(_05044_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11358_ (.I(_05044_),
    .Z(_00617_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11359_ (.I(_04959_),
    .Z(_05045_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11360_ (.I(_05045_),
    .Z(_05046_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11361_ (.I(_03864_),
    .Z(_05047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11362_ (.A1(_05047_),
    .A2(_05038_),
    .ZN(_05048_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11363_ (.I0(_05046_),
    .I1(\mod.u_cpu.rf_ram.memory[305][0] ),
    .S(_05048_),
    .Z(_05049_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11364_ (.I(_05049_),
    .Z(_00618_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11365_ (.I(_05031_),
    .Z(_05050_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11366_ (.I0(_05050_),
    .I1(\mod.u_cpu.rf_ram.memory[305][1] ),
    .S(_05048_),
    .Z(_05051_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11367_ (.I(_05051_),
    .Z(_00619_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11368_ (.A1(_04766_),
    .A2(_05038_),
    .ZN(_05052_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11369_ (.I0(_05046_),
    .I1(\mod.u_cpu.rf_ram.memory[304][0] ),
    .S(_05052_),
    .Z(_05053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11370_ (.I(_05053_),
    .Z(_00620_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11371_ (.I0(_05050_),
    .I1(\mod.u_cpu.rf_ram.memory[304][1] ),
    .S(_05052_),
    .Z(_05054_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11372_ (.I(_05054_),
    .Z(_00621_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11373_ (.A1(_04369_),
    .A2(_05020_),
    .ZN(_05055_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11374_ (.A1(_05022_),
    .A2(_05055_),
    .ZN(_05056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11375_ (.A1(_01968_),
    .A2(_05055_),
    .B(_05056_),
    .ZN(_00622_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11376_ (.I0(_05050_),
    .I1(\mod.u_cpu.rf_ram.memory[303][1] ),
    .S(_05055_),
    .Z(_05057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11377_ (.I(_05057_),
    .Z(_00623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11378_ (.I(_04995_),
    .Z(_05058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11379_ (.A1(_04775_),
    .A2(_05058_),
    .ZN(_05059_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11380_ (.I0(_05046_),
    .I1(\mod.u_cpu.rf_ram.memory[302][0] ),
    .S(_05059_),
    .Z(_05060_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11381_ (.I(_05060_),
    .Z(_00624_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11382_ (.I0(_05050_),
    .I1(\mod.u_cpu.rf_ram.memory[302][1] ),
    .S(_05059_),
    .Z(_05061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11383_ (.I(_05061_),
    .Z(_00625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11384_ (.A1(_03892_),
    .A2(_04779_),
    .ZN(_05062_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11385_ (.A1(_04377_),
    .A2(_05062_),
    .ZN(_05063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11386_ (.A1(_04817_),
    .A2(_05063_),
    .ZN(_05064_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11387_ (.A1(_01964_),
    .A2(_05063_),
    .B(_05064_),
    .ZN(_00626_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11388_ (.I(_04531_),
    .Z(_05065_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11389_ (.I0(\mod.u_cpu.rf_ram.memory[301][1] ),
    .I1(_05065_),
    .S(_05063_),
    .Z(_05066_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11390_ (.I(_05066_),
    .Z(_00627_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11391_ (.A1(_04784_),
    .A2(_05058_),
    .ZN(_05067_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11392_ (.I0(_05046_),
    .I1(\mod.u_cpu.rf_ram.memory[300][0] ),
    .S(_05067_),
    .Z(_05068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11393_ (.I(_05068_),
    .Z(_00628_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11394_ (.I(_05031_),
    .Z(_05069_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11395_ (.I0(_05069_),
    .I1(\mod.u_cpu.rf_ram.memory[300][1] ),
    .S(_05067_),
    .Z(_05070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11396_ (.I(_05070_),
    .Z(_00629_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11397_ (.I(_05045_),
    .Z(_05071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11398_ (.A1(_04196_),
    .A2(_03975_),
    .ZN(_05072_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11399_ (.I0(_05071_),
    .I1(\mod.u_cpu.rf_ram.memory[2][0] ),
    .S(_05072_),
    .Z(_05073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11400_ (.I(_05073_),
    .Z(_00630_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11401_ (.I0(_05069_),
    .I1(\mod.u_cpu.rf_ram.memory[2][1] ),
    .S(_05072_),
    .Z(_05074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11402_ (.I(_05074_),
    .Z(_00631_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11403_ (.A1(_04792_),
    .A2(_05058_),
    .ZN(_05075_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11404_ (.I0(_05071_),
    .I1(\mod.u_cpu.rf_ram.memory[298][0] ),
    .S(_05075_),
    .Z(_05076_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11405_ (.I(_05076_),
    .Z(_00632_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11406_ (.I0(_05069_),
    .I1(\mod.u_cpu.rf_ram.memory[298][1] ),
    .S(_05075_),
    .Z(_05077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11407_ (.I(_05077_),
    .Z(_00633_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11408_ (.I(_03712_),
    .Z(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11409_ (.A1(_05078_),
    .A2(_05062_),
    .ZN(_05079_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11410_ (.I0(\mod.u_cpu.rf_ram.memory[297][0] ),
    .I1(_04954_),
    .S(_05079_),
    .Z(_05080_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11411_ (.I(_05080_),
    .Z(_00634_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11412_ (.I0(\mod.u_cpu.rf_ram.memory[297][1] ),
    .I1(_05065_),
    .S(_05079_),
    .Z(_05081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11413_ (.I(_05081_),
    .Z(_00635_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11414_ (.A1(_04804_),
    .A2(_05058_),
    .ZN(_05082_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11415_ (.I0(_05071_),
    .I1(\mod.u_cpu.rf_ram.memory[296][0] ),
    .S(_05082_),
    .Z(_05083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11416_ (.I(_05083_),
    .Z(_00636_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11417_ (.I0(_05069_),
    .I1(\mod.u_cpu.rf_ram.memory[296][1] ),
    .S(_05082_),
    .Z(_05084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11418_ (.I(_05084_),
    .Z(_00637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11419_ (.A1(_04539_),
    .A2(_05020_),
    .ZN(_05085_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11420_ (.A1(_05022_),
    .A2(_05085_),
    .ZN(_05086_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11421_ (.A1(_01950_),
    .A2(_05085_),
    .B(_05086_),
    .ZN(_00638_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11422_ (.I(_05031_),
    .Z(_05087_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11423_ (.I0(_05087_),
    .I1(\mod.u_cpu.rf_ram.memory[295][1] ),
    .S(_05085_),
    .Z(_05088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11424_ (.I(_05088_),
    .Z(_00639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11425_ (.I(_04995_),
    .Z(_05089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11426_ (.A1(_04812_),
    .A2(_05089_),
    .ZN(_05090_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11427_ (.I0(_05071_),
    .I1(\mod.u_cpu.rf_ram.memory[294][0] ),
    .S(_05090_),
    .Z(_05091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11428_ (.I(_05091_),
    .Z(_00640_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11429_ (.I0(_05087_),
    .I1(\mod.u_cpu.rf_ram.memory[294][1] ),
    .S(_05090_),
    .Z(_05092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11430_ (.I(_05092_),
    .Z(_00641_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11431_ (.A1(_04412_),
    .A2(_05062_),
    .ZN(_05093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11432_ (.A1(_04817_),
    .A2(_05093_),
    .ZN(_05094_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11433_ (.A1(_01946_),
    .A2(_05093_),
    .B(_05094_),
    .ZN(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11434_ (.I0(\mod.u_cpu.rf_ram.memory[293][1] ),
    .I1(_05065_),
    .S(_05093_),
    .Z(_05095_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11435_ (.I(_05095_),
    .Z(_00643_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11436_ (.I(_05045_),
    .Z(_05096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11437_ (.A1(_04821_),
    .A2(_05089_),
    .ZN(_05097_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11438_ (.I0(_05096_),
    .I1(\mod.u_cpu.rf_ram.memory[292][0] ),
    .S(_05097_),
    .Z(_05098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11439_ (.I(_05098_),
    .Z(_00644_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11440_ (.I0(_05087_),
    .I1(\mod.u_cpu.rf_ram.memory[292][1] ),
    .S(_05097_),
    .Z(_05099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11441_ (.I(_05099_),
    .Z(_00645_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11442_ (.A1(_04965_),
    .A2(_05089_),
    .ZN(_05100_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11443_ (.I0(_05096_),
    .I1(\mod.u_cpu.rf_ram.memory[291][0] ),
    .S(_05100_),
    .Z(_05101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11444_ (.I(_05101_),
    .Z(_00646_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11445_ (.I0(_05087_),
    .I1(\mod.u_cpu.rf_ram.memory[291][1] ),
    .S(_05100_),
    .Z(_05102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11446_ (.I(_05102_),
    .Z(_00647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11447_ (.A1(_04831_),
    .A2(_05089_),
    .ZN(_05103_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11448_ (.I0(_05096_),
    .I1(\mod.u_cpu.rf_ram.memory[290][0] ),
    .S(_05103_),
    .Z(_05104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11449_ (.I(_05104_),
    .Z(_00648_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11450_ (.I(_03732_),
    .Z(_05105_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11451_ (.I(_05105_),
    .Z(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11452_ (.I(_05106_),
    .Z(_05107_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11453_ (.I(_05107_),
    .Z(_05108_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11454_ (.I0(_05108_),
    .I1(\mod.u_cpu.rf_ram.memory[290][1] ),
    .S(_05103_),
    .Z(_05109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11455_ (.I(_05109_),
    .Z(_00649_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11456_ (.I(_04195_),
    .Z(_05110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11457_ (.A1(_05110_),
    .A2(_03782_),
    .ZN(_05111_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11458_ (.I0(_05096_),
    .I1(\mod.u_cpu.rf_ram.memory[28][0] ),
    .S(_05111_),
    .Z(_05112_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11459_ (.I(_05112_),
    .Z(_00650_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11460_ (.I0(_05108_),
    .I1(\mod.u_cpu.rf_ram.memory[28][1] ),
    .S(_05111_),
    .Z(_05113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11461_ (.I(_05113_),
    .Z(_00651_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11462_ (.I(_05045_),
    .Z(_05114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11463_ (.A1(_04838_),
    .A2(_04996_),
    .ZN(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11464_ (.I0(_05114_),
    .I1(\mod.u_cpu.rf_ram.memory[288][0] ),
    .S(_05115_),
    .Z(_05116_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11465_ (.I(_05116_),
    .Z(_00652_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11466_ (.I0(_05108_),
    .I1(\mod.u_cpu.rf_ram.memory[288][1] ),
    .S(_05115_),
    .Z(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11467_ (.I(_05117_),
    .Z(_00653_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11468_ (.A1(_03993_),
    .A2(_04701_),
    .ZN(_05118_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11469_ (.I(_05118_),
    .Z(_05119_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11470_ (.I(_05119_),
    .Z(_05120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11471_ (.A1(_04700_),
    .A2(_05120_),
    .ZN(_05121_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11472_ (.A1(_05022_),
    .A2(_05121_),
    .ZN(_05122_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11473_ (.A1(_02002_),
    .A2(_05121_),
    .B(_05122_),
    .ZN(_00654_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11474_ (.I0(_05108_),
    .I1(\mod.u_cpu.rf_ram.memory[287][1] ),
    .S(_05121_),
    .Z(_05123_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11475_ (.I(_05123_),
    .Z(_00655_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11476_ (.I(_05118_),
    .Z(_05124_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11477_ (.I(_05124_),
    .Z(_05125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11478_ (.A1(_04852_),
    .A2(_05125_),
    .ZN(_05126_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11479_ (.I0(_05114_),
    .I1(\mod.u_cpu.rf_ram.memory[286][0] ),
    .S(_05126_),
    .Z(_05127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11480_ (.I(_05127_),
    .Z(_00656_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11481_ (.I(_05107_),
    .Z(_05128_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11482_ (.I0(_05128_),
    .I1(\mod.u_cpu.rf_ram.memory[286][1] ),
    .S(_05126_),
    .Z(_05129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11483_ (.I(_05129_),
    .Z(_00657_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11484_ (.I(_05119_),
    .Z(_05130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11485_ (.A1(_04994_),
    .A2(_05130_),
    .ZN(_05131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11486_ (.I(_03773_),
    .Z(_05132_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11487_ (.I(_05132_),
    .Z(_05133_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11488_ (.A1(_05133_),
    .A2(_05131_),
    .ZN(_05134_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11489_ (.A1(_01999_),
    .A2(_05131_),
    .B(_05134_),
    .ZN(_00658_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11490_ (.I0(_05128_),
    .I1(\mod.u_cpu.rf_ram.memory[285][1] ),
    .S(_05131_),
    .Z(_05135_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11491_ (.I(_05135_),
    .Z(_00659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11492_ (.A1(_04859_),
    .A2(_05125_),
    .ZN(_05136_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11493_ (.I0(_05114_),
    .I1(\mod.u_cpu.rf_ram.memory[284][0] ),
    .S(_05136_),
    .Z(_05137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11494_ (.I(_05137_),
    .Z(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11495_ (.I0(_05128_),
    .I1(\mod.u_cpu.rf_ram.memory[284][1] ),
    .S(_05136_),
    .Z(_05138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11496_ (.I(_05138_),
    .Z(_00661_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11497_ (.I(_03789_),
    .Z(_05139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11498_ (.A1(_05139_),
    .A2(_05125_),
    .ZN(_05140_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11499_ (.I0(_05114_),
    .I1(\mod.u_cpu.rf_ram.memory[283][0] ),
    .S(_05140_),
    .Z(_05141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11500_ (.I(_05141_),
    .Z(_00662_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11501_ (.I0(_05128_),
    .I1(\mod.u_cpu.rf_ram.memory[283][1] ),
    .S(_05140_),
    .Z(_05142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11502_ (.I(_05142_),
    .Z(_00663_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11503_ (.I(_04959_),
    .Z(_05143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11504_ (.I(_05143_),
    .Z(_05144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11505_ (.A1(_04868_),
    .A2(_05125_),
    .ZN(_05145_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11506_ (.I0(_05144_),
    .I1(\mod.u_cpu.rf_ram.memory[282][0] ),
    .S(_05145_),
    .Z(_05146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11507_ (.I(_05146_),
    .Z(_00664_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11508_ (.I(_05107_),
    .Z(_05147_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11509_ (.I0(_05147_),
    .I1(\mod.u_cpu.rf_ram.memory[282][1] ),
    .S(_05145_),
    .Z(_05148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11510_ (.I(_05148_),
    .Z(_00665_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11511_ (.I(_05124_),
    .Z(_05149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11512_ (.A1(_04873_),
    .A2(_05149_),
    .ZN(_05150_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11513_ (.I0(_05144_),
    .I1(\mod.u_cpu.rf_ram.memory[281][0] ),
    .S(_05150_),
    .Z(_05151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11514_ (.I(_05151_),
    .Z(_00666_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11515_ (.I0(_05147_),
    .I1(\mod.u_cpu.rf_ram.memory[281][1] ),
    .S(_05150_),
    .Z(_05152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11516_ (.I(_05152_),
    .Z(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11517_ (.A1(_04732_),
    .A2(_05149_),
    .ZN(_05153_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11518_ (.I0(_05144_),
    .I1(\mod.u_cpu.rf_ram.memory[280][0] ),
    .S(_05153_),
    .Z(_05154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11519_ (.I(_05154_),
    .Z(_00668_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11520_ (.I0(_05147_),
    .I1(\mod.u_cpu.rf_ram.memory[280][1] ),
    .S(_05153_),
    .Z(_05155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11521_ (.I(_05155_),
    .Z(_00669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11522_ (.A1(_05110_),
    .A2(_03791_),
    .ZN(_05156_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11523_ (.I0(_05144_),
    .I1(\mod.u_cpu.rf_ram.memory[27][0] ),
    .S(_05156_),
    .Z(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11524_ (.I(_05157_),
    .Z(_00670_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11525_ (.I0(_05147_),
    .I1(\mod.u_cpu.rf_ram.memory[27][1] ),
    .S(_05156_),
    .Z(_05158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11526_ (.I(_05158_),
    .Z(_00671_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11527_ (.I(_05143_),
    .Z(_05159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11528_ (.A1(_04741_),
    .A2(_05149_),
    .ZN(_05160_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11529_ (.I0(_05159_),
    .I1(\mod.u_cpu.rf_ram.memory[278][0] ),
    .S(_05160_),
    .Z(_05161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11530_ (.I(_05161_),
    .Z(_00672_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11531_ (.I(_05107_),
    .Z(_05162_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11532_ (.I0(_05162_),
    .I1(\mod.u_cpu.rf_ram.memory[278][1] ),
    .S(_05160_),
    .Z(_05163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11533_ (.I(_05163_),
    .Z(_00673_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11534_ (.I(_03835_),
    .Z(_05164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11535_ (.A1(_05164_),
    .A2(_05130_),
    .ZN(_05165_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11536_ (.A1(_05133_),
    .A2(_05165_),
    .ZN(_05166_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11537_ (.A1(_01982_),
    .A2(_05165_),
    .B(_05166_),
    .ZN(_00674_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11538_ (.I0(_05162_),
    .I1(\mod.u_cpu.rf_ram.memory[277][1] ),
    .S(_05165_),
    .Z(_05167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11539_ (.I(_05167_),
    .Z(_00675_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11540_ (.A1(_04749_),
    .A2(_05149_),
    .ZN(_05168_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11541_ (.I0(_05159_),
    .I1(\mod.u_cpu.rf_ram.memory[276][0] ),
    .S(_05168_),
    .Z(_05169_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11542_ (.I(_05169_),
    .Z(_00676_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11543_ (.I0(_05162_),
    .I1(\mod.u_cpu.rf_ram.memory[276][1] ),
    .S(_05168_),
    .Z(_05170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11544_ (.I(_05170_),
    .Z(_00677_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11545_ (.I(_05124_),
    .Z(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11546_ (.A1(_05037_),
    .A2(_05171_),
    .ZN(_05172_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11547_ (.I0(_05159_),
    .I1(\mod.u_cpu.rf_ram.memory[275][0] ),
    .S(_05172_),
    .Z(_05173_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11548_ (.I(_05173_),
    .Z(_00678_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11549_ (.I0(_05162_),
    .I1(\mod.u_cpu.rf_ram.memory[275][1] ),
    .S(_05172_),
    .Z(_05174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11550_ (.I(_05174_),
    .Z(_00679_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11551_ (.A1(_04758_),
    .A2(_05171_),
    .ZN(_05175_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11552_ (.I0(_05159_),
    .I1(\mod.u_cpu.rf_ram.memory[274][0] ),
    .S(_05175_),
    .Z(_05176_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11553_ (.I(_05176_),
    .Z(_00680_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11554_ (.I(_05106_),
    .Z(_05177_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11555_ (.I(_05177_),
    .Z(_05178_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11556_ (.I0(_05178_),
    .I1(\mod.u_cpu.rf_ram.memory[274][1] ),
    .S(_05175_),
    .Z(_05179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11557_ (.I(_05179_),
    .Z(_00681_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11558_ (.I(_05143_),
    .Z(_05180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11559_ (.A1(_05047_),
    .A2(_05171_),
    .ZN(_05181_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11560_ (.I0(_05180_),
    .I1(\mod.u_cpu.rf_ram.memory[273][0] ),
    .S(_05181_),
    .Z(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11561_ (.I(_05182_),
    .Z(_00682_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11562_ (.I0(_05178_),
    .I1(\mod.u_cpu.rf_ram.memory[273][1] ),
    .S(_05181_),
    .Z(_05183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11563_ (.I(_05183_),
    .Z(_00683_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11564_ (.A1(_04766_),
    .A2(_05171_),
    .ZN(_05184_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11565_ (.I0(_05180_),
    .I1(\mod.u_cpu.rf_ram.memory[272][0] ),
    .S(_05184_),
    .Z(_05185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11566_ (.I(_05185_),
    .Z(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11567_ (.I0(_05178_),
    .I1(\mod.u_cpu.rf_ram.memory[272][1] ),
    .S(_05184_),
    .Z(_05186_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11568_ (.I(_05186_),
    .Z(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11569_ (.I(_04066_),
    .Z(_05187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11570_ (.A1(_05187_),
    .A2(_05130_),
    .ZN(_05188_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11571_ (.A1(_05133_),
    .A2(_05188_),
    .ZN(_05189_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11572_ (.A1(_02028_),
    .A2(_05188_),
    .B(_05189_),
    .ZN(_00686_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11573_ (.I0(_05178_),
    .I1(\mod.u_cpu.rf_ram.memory[271][1] ),
    .S(_05188_),
    .Z(_05190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11574_ (.I(_05190_),
    .Z(_00687_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11575_ (.I(_05119_),
    .Z(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11576_ (.A1(_04775_),
    .A2(_05191_),
    .ZN(_05192_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11577_ (.I0(_05180_),
    .I1(\mod.u_cpu.rf_ram.memory[270][0] ),
    .S(_05192_),
    .Z(_05193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11578_ (.I(_05193_),
    .Z(_00688_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11579_ (.I(_05177_),
    .Z(_05194_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11580_ (.I0(_05194_),
    .I1(\mod.u_cpu.rf_ram.memory[270][1] ),
    .S(_05192_),
    .Z(_05195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11581_ (.I(_05195_),
    .Z(_00689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11582_ (.A1(_05110_),
    .A2(_03797_),
    .ZN(_05196_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11583_ (.I0(_05180_),
    .I1(\mod.u_cpu.rf_ram.memory[26][0] ),
    .S(_05196_),
    .Z(_05197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11584_ (.I(_05197_),
    .Z(_00690_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11585_ (.I0(_05194_),
    .I1(\mod.u_cpu.rf_ram.memory[26][1] ),
    .S(_05196_),
    .Z(_05198_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11586_ (.I(_05198_),
    .Z(_00691_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11587_ (.I(_05143_),
    .Z(_05199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11588_ (.A1(_04784_),
    .A2(_05191_),
    .ZN(_05200_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11589_ (.I0(_05199_),
    .I1(\mod.u_cpu.rf_ram.memory[268][0] ),
    .S(_05200_),
    .Z(_05201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11590_ (.I(_05201_),
    .Z(_00692_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11591_ (.I0(_05194_),
    .I1(\mod.u_cpu.rf_ram.memory[268][1] ),
    .S(_05200_),
    .Z(_05202_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11592_ (.I(_05202_),
    .Z(_00693_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11593_ (.A1(_04930_),
    .A2(_05191_),
    .ZN(_05203_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11594_ (.I0(_05199_),
    .I1(\mod.u_cpu.rf_ram.memory[267][0] ),
    .S(_05203_),
    .Z(_05204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11595_ (.I(_05204_),
    .Z(_00694_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11596_ (.I0(_05194_),
    .I1(\mod.u_cpu.rf_ram.memory[267][1] ),
    .S(_05203_),
    .Z(_05205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11597_ (.I(_05205_),
    .Z(_00695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11598_ (.A1(_04792_),
    .A2(_05191_),
    .ZN(_05206_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11599_ (.I0(_05199_),
    .I1(\mod.u_cpu.rf_ram.memory[266][0] ),
    .S(_05206_),
    .Z(_05207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11600_ (.I(_05207_),
    .Z(_00696_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11601_ (.I(_05177_),
    .Z(_05208_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11602_ (.I0(_05208_),
    .I1(\mod.u_cpu.rf_ram.memory[266][1] ),
    .S(_05206_),
    .Z(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11603_ (.I(_05209_),
    .Z(_00697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11604_ (.A1(_03723_),
    .A2(_04779_),
    .ZN(_05210_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11605_ (.A1(_05078_),
    .A2(_05210_),
    .ZN(_05211_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11606_ (.I0(\mod.u_cpu.rf_ram.memory[265][0] ),
    .I1(_04954_),
    .S(_05211_),
    .Z(_05212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11607_ (.I(_05212_),
    .Z(_00698_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11608_ (.I0(\mod.u_cpu.rf_ram.memory[265][1] ),
    .I1(_05065_),
    .S(_05211_),
    .Z(_05213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11609_ (.I(_05213_),
    .Z(_00699_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11610_ (.I(_05119_),
    .Z(_05214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11611_ (.A1(_04804_),
    .A2(_05214_),
    .ZN(_05215_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11612_ (.I0(_05199_),
    .I1(\mod.u_cpu.rf_ram.memory[264][0] ),
    .S(_05215_),
    .Z(_05216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11613_ (.I(_05216_),
    .Z(_00700_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11614_ (.I0(_05208_),
    .I1(\mod.u_cpu.rf_ram.memory[264][1] ),
    .S(_05215_),
    .Z(_05217_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11615_ (.I(_05217_),
    .Z(_00701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11616_ (.A1(_04539_),
    .A2(_05130_),
    .ZN(_05218_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11617_ (.A1(_05133_),
    .A2(_05218_),
    .ZN(_05219_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11618_ (.A1(_02015_),
    .A2(_05218_),
    .B(_05219_),
    .ZN(_00702_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11619_ (.I0(_05208_),
    .I1(\mod.u_cpu.rf_ram.memory[263][1] ),
    .S(_05218_),
    .Z(_05220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11620_ (.I(_05220_),
    .Z(_00703_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11621_ (.I(_04959_),
    .Z(_05221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11622_ (.I(_05221_),
    .Z(_05222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11623_ (.A1(_04812_),
    .A2(_05214_),
    .ZN(_05223_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11624_ (.I0(_05222_),
    .I1(\mod.u_cpu.rf_ram.memory[262][0] ),
    .S(_05223_),
    .Z(_05224_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11625_ (.I(_05224_),
    .Z(_00704_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11626_ (.I0(_05208_),
    .I1(\mod.u_cpu.rf_ram.memory[262][1] ),
    .S(_05223_),
    .Z(_05225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11627_ (.I(_05225_),
    .Z(_00705_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11628_ (.I(_04106_),
    .Z(_05226_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11629_ (.A1(_05226_),
    .A2(_05210_),
    .ZN(_05227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11630_ (.A1(_04817_),
    .A2(_05227_),
    .ZN(_05228_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11631_ (.A1(_02012_),
    .A2(_05227_),
    .B(_05228_),
    .ZN(_00706_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11632_ (.I(_03733_),
    .Z(_05229_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11633_ (.I(_05229_),
    .Z(_05230_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11634_ (.I0(\mod.u_cpu.rf_ram.memory[261][1] ),
    .I1(_05230_),
    .S(_05227_),
    .Z(_05231_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11635_ (.I(_05231_),
    .Z(_00707_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11636_ (.A1(_04821_),
    .A2(_05214_),
    .ZN(_05232_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11637_ (.I0(_05222_),
    .I1(\mod.u_cpu.rf_ram.memory[260][0] ),
    .S(_05232_),
    .Z(_05233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11638_ (.I(_05233_),
    .Z(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11639_ (.I(_05177_),
    .Z(_05234_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11640_ (.I0(_05234_),
    .I1(\mod.u_cpu.rf_ram.memory[260][1] ),
    .S(_05232_),
    .Z(_05235_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11641_ (.I(_05235_),
    .Z(_00709_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11642_ (.A1(_05110_),
    .A2(_04026_),
    .ZN(_05236_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11643_ (.I0(_05222_),
    .I1(\mod.u_cpu.rf_ram.memory[25][0] ),
    .S(_05236_),
    .Z(_05237_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11644_ (.I(_05237_),
    .Z(_00710_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11645_ (.I0(_05234_),
    .I1(\mod.u_cpu.rf_ram.memory[25][1] ),
    .S(_05236_),
    .Z(_05238_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11646_ (.I(_05238_),
    .Z(_00711_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11647_ (.I(_04195_),
    .Z(_05239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11648_ (.A1(_05239_),
    .A2(_03805_),
    .ZN(_05240_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11649_ (.I0(_05222_),
    .I1(\mod.u_cpu.rf_ram.memory[24][0] ),
    .S(_05240_),
    .Z(_05241_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11650_ (.I(_05241_),
    .Z(_00712_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11651_ (.I0(_05234_),
    .I1(\mod.u_cpu.rf_ram.memory[24][1] ),
    .S(_05240_),
    .Z(_05242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11652_ (.I(_05242_),
    .Z(_00713_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11653_ (.I(_05221_),
    .Z(_05243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11654_ (.A1(_04831_),
    .A2(_05214_),
    .ZN(_05244_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11655_ (.I0(_05243_),
    .I1(\mod.u_cpu.rf_ram.memory[258][0] ),
    .S(_05244_),
    .Z(_05245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11656_ (.I(_05245_),
    .Z(_00714_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11657_ (.I0(_05234_),
    .I1(\mod.u_cpu.rf_ram.memory[258][1] ),
    .S(_05244_),
    .Z(_05246_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11658_ (.I(_05246_),
    .Z(_00715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11659_ (.A1(_04973_),
    .A2(_05120_),
    .ZN(_05247_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11660_ (.I0(_05243_),
    .I1(\mod.u_cpu.rf_ram.memory[257][0] ),
    .S(_05247_),
    .Z(_05248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11661_ (.I(_05248_),
    .Z(_00716_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11662_ (.I(_05106_),
    .Z(_05249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11663_ (.I(_05249_),
    .Z(_05250_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11664_ (.I0(_05250_),
    .I1(\mod.u_cpu.rf_ram.memory[257][1] ),
    .S(_05247_),
    .Z(_05251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11665_ (.I(_05251_),
    .Z(_00717_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11666_ (.A1(_03665_),
    .A2(_04224_),
    .ZN(_05252_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11667_ (.A1(_04226_),
    .A2(_05252_),
    .Z(_05253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11668_ (.I(_05253_),
    .Z(_05254_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11669_ (.I(_05254_),
    .Z(_05255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11670_ (.A1(_04868_),
    .A2(_05255_),
    .ZN(_05256_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11671_ (.I0(_05243_),
    .I1(\mod.u_cpu.rf_ram.memory[250][0] ),
    .S(_05256_),
    .Z(_05257_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11672_ (.I(_05257_),
    .Z(_00718_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11673_ (.I0(_05250_),
    .I1(\mod.u_cpu.rf_ram.memory[250][1] ),
    .S(_05256_),
    .Z(_05258_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11674_ (.I(_05258_),
    .Z(_00719_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11675_ (.A1(_04838_),
    .A2(_05120_),
    .ZN(_05259_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11676_ (.I0(_05243_),
    .I1(\mod.u_cpu.rf_ram.memory[256][0] ),
    .S(_05259_),
    .Z(_05260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11677_ (.I(_05260_),
    .Z(_00720_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11678_ (.I0(_05250_),
    .I1(\mod.u_cpu.rf_ram.memory[256][1] ),
    .S(_05259_),
    .Z(_05261_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11679_ (.I(_05261_),
    .Z(_00721_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11680_ (.I(_05253_),
    .Z(_05262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11681_ (.I(_05262_),
    .Z(_05263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11682_ (.A1(_04700_),
    .A2(_05263_),
    .ZN(_05264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11683_ (.I(_05132_),
    .Z(_05265_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11684_ (.A1(_05265_),
    .A2(_05264_),
    .ZN(_05266_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11685_ (.A1(_02273_),
    .A2(_05264_),
    .B(_05266_),
    .ZN(_00722_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11686_ (.I0(_05250_),
    .I1(\mod.u_cpu.rf_ram.memory[255][1] ),
    .S(_05264_),
    .Z(_05267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11687_ (.I(_05267_),
    .Z(_00723_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11688_ (.I(_05221_),
    .Z(_05268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11689_ (.A1(_05139_),
    .A2(_05255_),
    .ZN(_05269_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11690_ (.I0(_05268_),
    .I1(\mod.u_cpu.rf_ram.memory[251][0] ),
    .S(_05269_),
    .Z(_05270_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11691_ (.I(_05270_),
    .Z(_00724_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11692_ (.I(_05249_),
    .Z(_05271_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11693_ (.I0(_05271_),
    .I1(\mod.u_cpu.rf_ram.memory[251][1] ),
    .S(_05269_),
    .Z(_05272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11694_ (.I(_05272_),
    .Z(_00725_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11695_ (.A1(_04852_),
    .A2(_05255_),
    .ZN(_05273_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11696_ (.I0(_05268_),
    .I1(\mod.u_cpu.rf_ram.memory[254][0] ),
    .S(_05273_),
    .Z(_05274_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11697_ (.I(_05274_),
    .Z(_00726_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11698_ (.I0(_05271_),
    .I1(\mod.u_cpu.rf_ram.memory[254][1] ),
    .S(_05273_),
    .Z(_05275_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11699_ (.I(_05275_),
    .Z(_00727_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11700_ (.A1(_04859_),
    .A2(_05255_),
    .ZN(_05276_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11701_ (.I0(_05268_),
    .I1(\mod.u_cpu.rf_ram.memory[252][0] ),
    .S(_05276_),
    .Z(_05277_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11702_ (.I(_05277_),
    .Z(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11703_ (.I0(_05271_),
    .I1(\mod.u_cpu.rf_ram.memory[252][1] ),
    .S(_05276_),
    .Z(_05278_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11704_ (.I(_05278_),
    .Z(_00729_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11705_ (.I(_05262_),
    .Z(_05279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11706_ (.A1(_04994_),
    .A2(_05279_),
    .ZN(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11707_ (.A1(_05265_),
    .A2(_05280_),
    .ZN(_05281_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11708_ (.A1(_02269_),
    .A2(_05280_),
    .B(_05281_),
    .ZN(_00730_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11709_ (.I0(_05271_),
    .I1(\mod.u_cpu.rf_ram.memory[253][1] ),
    .S(_05280_),
    .Z(_05282_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11710_ (.I(_05282_),
    .Z(_00731_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11711_ (.I(_03803_),
    .Z(_05283_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11712_ (.I(_05254_),
    .Z(_05284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11713_ (.A1(_05283_),
    .A2(_05284_),
    .ZN(_05285_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11714_ (.I0(_05268_),
    .I1(\mod.u_cpu.rf_ram.memory[248][0] ),
    .S(_05285_),
    .Z(_05286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11715_ (.I(_05286_),
    .Z(_00732_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11716_ (.I(_05249_),
    .Z(_05287_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11717_ (.I0(_05287_),
    .I1(\mod.u_cpu.rf_ram.memory[248][1] ),
    .S(_05285_),
    .Z(_05288_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11718_ (.I(_05288_),
    .Z(_00733_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11719_ (.I(_05221_),
    .Z(_05289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11720_ (.A1(_05037_),
    .A2(_05284_),
    .ZN(_05290_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11721_ (.I0(_05289_),
    .I1(\mod.u_cpu.rf_ram.memory[243][0] ),
    .S(_05290_),
    .Z(_05291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11722_ (.I(_05291_),
    .Z(_00734_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11723_ (.I0(_05287_),
    .I1(\mod.u_cpu.rf_ram.memory[243][1] ),
    .S(_05290_),
    .Z(_05292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11724_ (.I(_05292_),
    .Z(_00735_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11725_ (.I(_03857_),
    .Z(_05293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11726_ (.A1(_05293_),
    .A2(_05284_),
    .ZN(_05294_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11727_ (.I0(_05289_),
    .I1(\mod.u_cpu.rf_ram.memory[242][0] ),
    .S(_05294_),
    .Z(_05295_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11728_ (.I(_05295_),
    .Z(_00736_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11729_ (.I0(_05287_),
    .I1(\mod.u_cpu.rf_ram.memory[242][1] ),
    .S(_05294_),
    .Z(_05296_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11730_ (.I(_05296_),
    .Z(_00737_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11731_ (.A1(_05047_),
    .A2(_05284_),
    .ZN(_05297_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11732_ (.I0(_05289_),
    .I1(\mod.u_cpu.rf_ram.memory[241][0] ),
    .S(_05297_),
    .Z(_05298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11733_ (.I(_05298_),
    .Z(_00738_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11734_ (.I0(_05287_),
    .I1(\mod.u_cpu.rf_ram.memory[241][1] ),
    .S(_05297_),
    .Z(_05299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11735_ (.I(_05299_),
    .Z(_00739_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11736_ (.I(_03871_),
    .Z(_05300_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11737_ (.I(_05254_),
    .Z(_05301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11738_ (.A1(_05300_),
    .A2(_05301_),
    .ZN(_05302_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11739_ (.I0(_05289_),
    .I1(\mod.u_cpu.rf_ram.memory[240][0] ),
    .S(_05302_),
    .Z(_05303_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11740_ (.I(_05303_),
    .Z(_00740_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11741_ (.I(_05249_),
    .Z(_05304_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11742_ (.I0(_05304_),
    .I1(\mod.u_cpu.rf_ram.memory[240][1] ),
    .S(_05302_),
    .Z(_05305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11743_ (.I(_05305_),
    .Z(_00741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11744_ (.A1(_04983_),
    .A2(_03823_),
    .ZN(_05306_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11745_ (.A1(_05265_),
    .A2(_05306_),
    .ZN(_05307_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11746_ (.A1(_02412_),
    .A2(_05306_),
    .B(_05307_),
    .ZN(_00742_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11747_ (.I0(_05304_),
    .I1(\mod.u_cpu.rf_ram.memory[23][1] ),
    .S(_05306_),
    .Z(_05308_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11748_ (.I(_05308_),
    .Z(_00743_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11749_ (.I(_03696_),
    .Z(_05309_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11750_ (.I(_05309_),
    .Z(_05310_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11751_ (.I(_05310_),
    .Z(_05311_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11752_ (.I(_03884_),
    .Z(_05312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11753_ (.A1(_05312_),
    .A2(_05301_),
    .ZN(_05313_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11754_ (.I0(_05311_),
    .I1(\mod.u_cpu.rf_ram.memory[238][0] ),
    .S(_05313_),
    .Z(_05314_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11755_ (.I(_05314_),
    .Z(_00744_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11756_ (.I0(_05304_),
    .I1(\mod.u_cpu.rf_ram.memory[238][1] ),
    .S(_05313_),
    .Z(_05315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11757_ (.I(_05315_),
    .Z(_00745_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11758_ (.A1(_05187_),
    .A2(_05279_),
    .ZN(_05316_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11759_ (.A1(_05265_),
    .A2(_05316_),
    .ZN(_05317_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11760_ (.A1(_02250_),
    .A2(_05316_),
    .B(_05317_),
    .ZN(_00746_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11761_ (.I0(_05304_),
    .I1(\mod.u_cpu.rf_ram.memory[239][1] ),
    .S(_05316_),
    .Z(_05318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11762_ (.I(_05318_),
    .Z(_00747_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11763_ (.I(_05252_),
    .Z(_05319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11764_ (.A1(_04227_),
    .A2(_05319_),
    .ZN(_05320_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11765_ (.A1(_04377_),
    .A2(_05320_),
    .ZN(_05321_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11766_ (.I(_03944_),
    .Z(_05322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11767_ (.A1(_05322_),
    .A2(_05321_),
    .ZN(_05323_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11768_ (.A1(_02246_),
    .A2(_05321_),
    .B(_05323_),
    .ZN(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11769_ (.I0(\mod.u_cpu.rf_ram.memory[237][1] ),
    .I1(_05230_),
    .S(_05321_),
    .Z(_05324_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11770_ (.I(_05324_),
    .Z(_00749_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11771_ (.I(_03903_),
    .Z(_05325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11772_ (.A1(_05325_),
    .A2(_05301_),
    .ZN(_05326_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11773_ (.I0(_05311_),
    .I1(\mod.u_cpu.rf_ram.memory[236][0] ),
    .S(_05326_),
    .Z(_05327_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11774_ (.I(_05327_),
    .Z(_00750_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11775_ (.I(_05106_),
    .Z(_05328_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11776_ (.I(_05328_),
    .Z(_05329_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11777_ (.I0(_05329_),
    .I1(\mod.u_cpu.rf_ram.memory[236][1] ),
    .S(_05326_),
    .Z(_05330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11778_ (.I(_05330_),
    .Z(_00751_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11779_ (.A1(_04930_),
    .A2(_05301_),
    .ZN(_05331_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11780_ (.I0(_05311_),
    .I1(\mod.u_cpu.rf_ram.memory[235][0] ),
    .S(_05331_),
    .Z(_05332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11781_ (.I(_05332_),
    .Z(_00752_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11782_ (.I0(_05329_),
    .I1(\mod.u_cpu.rf_ram.memory[235][1] ),
    .S(_05331_),
    .Z(_05333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11783_ (.I(_05333_),
    .Z(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11784_ (.I(_03917_),
    .Z(_05334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11785_ (.I(_05262_),
    .Z(_05335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11786_ (.A1(_05334_),
    .A2(_05335_),
    .ZN(_05336_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11787_ (.I0(_05311_),
    .I1(\mod.u_cpu.rf_ram.memory[234][0] ),
    .S(_05336_),
    .Z(_05337_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11788_ (.I(_05337_),
    .Z(_00754_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11789_ (.I0(_05329_),
    .I1(\mod.u_cpu.rf_ram.memory[234][1] ),
    .S(_05336_),
    .Z(_05338_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11790_ (.I(_05338_),
    .Z(_00755_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11791_ (.A1(_05078_),
    .A2(_05320_),
    .ZN(_05339_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11792_ (.I0(\mod.u_cpu.rf_ram.memory[233][0] ),
    .I1(_04954_),
    .S(_05339_),
    .Z(_05340_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11793_ (.I(_05340_),
    .Z(_00756_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11794_ (.I0(\mod.u_cpu.rf_ram.memory[233][1] ),
    .I1(_05230_),
    .S(_05339_),
    .Z(_05341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11795_ (.I(_05341_),
    .Z(_00757_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11796_ (.I(_05310_),
    .Z(_05342_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11797_ (.I(_03931_),
    .Z(_05343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11798_ (.A1(_05343_),
    .A2(_05335_),
    .ZN(_05344_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11799_ (.I0(_05342_),
    .I1(\mod.u_cpu.rf_ram.memory[232][0] ),
    .S(_05344_),
    .Z(_05345_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11800_ (.I(_05345_),
    .Z(_00758_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11801_ (.I0(_05329_),
    .I1(\mod.u_cpu.rf_ram.memory[232][1] ),
    .S(_05344_),
    .Z(_05346_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11802_ (.I(_05346_),
    .Z(_00759_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11803_ (.A1(_04539_),
    .A2(_05279_),
    .ZN(_05347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11804_ (.I(_05132_),
    .Z(_05348_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11805_ (.A1(_05348_),
    .A2(_05347_),
    .ZN(_05349_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11806_ (.A1(_02237_),
    .A2(_05347_),
    .B(_05349_),
    .ZN(_00760_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11807_ (.I(_05328_),
    .Z(_05350_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11808_ (.I0(_05350_),
    .I1(\mod.u_cpu.rf_ram.memory[231][1] ),
    .S(_05347_),
    .Z(_05351_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11809_ (.I(_05351_),
    .Z(_00761_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11810_ (.A1(_04808_),
    .A2(_03866_),
    .ZN(_05352_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11811_ (.I0(_05342_),
    .I1(\mod.u_cpu.rf_ram.memory[49][0] ),
    .S(_05352_),
    .Z(_05353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11812_ (.I(_05353_),
    .Z(_00762_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11813_ (.I0(_05350_),
    .I1(\mod.u_cpu.rf_ram.memory[49][1] ),
    .S(_05352_),
    .Z(_05354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11814_ (.I(_05354_),
    .Z(_00763_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11815_ (.I(_03949_),
    .Z(_05355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11816_ (.A1(_05355_),
    .A2(_05335_),
    .ZN(_05356_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11817_ (.I0(_05342_),
    .I1(\mod.u_cpu.rf_ram.memory[230][0] ),
    .S(_05356_),
    .Z(_05357_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11818_ (.I(_05357_),
    .Z(_00764_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11819_ (.I0(_05350_),
    .I1(\mod.u_cpu.rf_ram.memory[230][1] ),
    .S(_05356_),
    .Z(_05358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11820_ (.I(_05358_),
    .Z(_00765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11821_ (.A1(_05239_),
    .A2(_03829_),
    .ZN(_05359_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11822_ (.I0(_05342_),
    .I1(\mod.u_cpu.rf_ram.memory[22][0] ),
    .S(_05359_),
    .Z(_05360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11823_ (.I(_05360_),
    .Z(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11824_ (.I0(_05350_),
    .I1(\mod.u_cpu.rf_ram.memory[22][1] ),
    .S(_05359_),
    .Z(_05361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11825_ (.I(_05361_),
    .Z(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11826_ (.A1(_04294_),
    .A2(_03942_),
    .ZN(_05362_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11827_ (.A1(_05348_),
    .A2(_05362_),
    .ZN(_05363_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11828_ (.A1(_02430_),
    .A2(_05362_),
    .B(_05363_),
    .ZN(_00768_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11829_ (.I(_05328_),
    .Z(_05364_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11830_ (.I0(_05364_),
    .I1(\mod.u_cpu.rf_ram.memory[39][1] ),
    .S(_05362_),
    .Z(_05365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11831_ (.I(_05365_),
    .Z(_00769_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11832_ (.I(_05310_),
    .Z(_05366_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11833_ (.I(_03959_),
    .Z(_05367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11834_ (.A1(_05367_),
    .A2(_05335_),
    .ZN(_05368_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11835_ (.I0(_05366_),
    .I1(\mod.u_cpu.rf_ram.memory[228][0] ),
    .S(_05368_),
    .Z(_05369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11836_ (.I(_05369_),
    .Z(_00770_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11837_ (.I0(_05364_),
    .I1(\mod.u_cpu.rf_ram.memory[228][1] ),
    .S(_05368_),
    .Z(_05370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11838_ (.I(_05370_),
    .Z(_00771_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11839_ (.A1(_03662_),
    .A2(_04223_),
    .A3(_03753_),
    .ZN(_05371_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11840_ (.A1(_03993_),
    .A2(_05371_),
    .ZN(_05372_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11841_ (.I(_05372_),
    .Z(_05373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11842_ (.I(_05373_),
    .Z(_05374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11843_ (.A1(_04845_),
    .A2(_05374_),
    .ZN(_05375_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11844_ (.I0(_05366_),
    .I1(\mod.u_cpu.rf_ram.memory[159][0] ),
    .S(_05375_),
    .Z(_05376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11845_ (.I(_05376_),
    .Z(_00772_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11846_ (.I0(_05364_),
    .I1(\mod.u_cpu.rf_ram.memory[159][1] ),
    .S(_05375_),
    .Z(_05377_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11847_ (.I(_05377_),
    .Z(_00773_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11848_ (.A1(_04014_),
    .A2(_05374_),
    .ZN(_05378_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11849_ (.I0(_05366_),
    .I1(\mod.u_cpu.rf_ram.memory[149][0] ),
    .S(_05378_),
    .Z(_05379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11850_ (.I(_05379_),
    .Z(_00774_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11851_ (.I0(_05364_),
    .I1(\mod.u_cpu.rf_ram.memory[149][1] ),
    .S(_05378_),
    .Z(_05380_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11852_ (.I(_05380_),
    .Z(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11853_ (.A1(_05239_),
    .A2(_03951_),
    .ZN(_05381_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11854_ (.I0(_05366_),
    .I1(\mod.u_cpu.rf_ram.memory[6][0] ),
    .S(_05381_),
    .Z(_05382_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11855_ (.I(_05382_),
    .Z(_00776_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11856_ (.I(_05328_),
    .Z(_05383_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11857_ (.I0(_05383_),
    .I1(\mod.u_cpu.rf_ram.memory[6][1] ),
    .S(_05381_),
    .Z(_05384_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11858_ (.I(_05384_),
    .Z(_00777_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11859_ (.I(_05310_),
    .Z(_05385_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11860_ (.A1(_03726_),
    .A2(_04378_),
    .Z(_05386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11861_ (.I(_05386_),
    .Z(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11862_ (.I(_05387_),
    .Z(_05388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11863_ (.A1(_05355_),
    .A2(_05388_),
    .ZN(_05389_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11864_ (.I0(_05385_),
    .I1(\mod.u_cpu.rf_ram.memory[70][0] ),
    .S(_05389_),
    .Z(_05390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11865_ (.I(_05390_),
    .Z(_00778_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11866_ (.I0(_05383_),
    .I1(\mod.u_cpu.rf_ram.memory[70][1] ),
    .S(_05389_),
    .Z(_05391_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11867_ (.I(_05391_),
    .Z(_00779_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11868_ (.A1(_05343_),
    .A2(_05388_),
    .ZN(_05392_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11869_ (.I0(_05385_),
    .I1(\mod.u_cpu.rf_ram.memory[72][0] ),
    .S(_05392_),
    .Z(_05393_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11870_ (.I(_05393_),
    .Z(_00780_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11871_ (.I0(_05383_),
    .I1(\mod.u_cpu.rf_ram.memory[72][1] ),
    .S(_05392_),
    .Z(_05394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11872_ (.I(_05394_),
    .Z(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11873_ (.I(_03940_),
    .Z(_05395_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11874_ (.I(_05386_),
    .Z(_05396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11875_ (.I(_05396_),
    .Z(_05397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11876_ (.A1(_05395_),
    .A2(_05397_),
    .ZN(_05398_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11877_ (.A1(_05348_),
    .A2(_05398_),
    .ZN(_05399_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11878_ (.A1(_02357_),
    .A2(_05398_),
    .B(_05399_),
    .ZN(_00782_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11879_ (.I0(_05383_),
    .I1(\mod.u_cpu.rf_ram.memory[71][1] ),
    .S(_05398_),
    .Z(_05400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11880_ (.I(_05400_),
    .Z(_00783_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11881_ (.I(_05262_),
    .Z(_05401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11882_ (.A1(_04965_),
    .A2(_05401_),
    .ZN(_05402_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11883_ (.I0(_05385_),
    .I1(\mod.u_cpu.rf_ram.memory[227][0] ),
    .S(_05402_),
    .Z(_05403_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11884_ (.I(_05403_),
    .Z(_00784_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11885_ (.I(_05105_),
    .Z(_05404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11886_ (.I(_05404_),
    .Z(_05405_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11887_ (.I(_05405_),
    .Z(_05406_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11888_ (.I0(_05406_),
    .I1(\mod.u_cpu.rf_ram.memory[227][1] ),
    .S(_05402_),
    .Z(_05407_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11889_ (.I(_05407_),
    .Z(_00785_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11890_ (.I(_03973_),
    .Z(_05408_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11891_ (.A1(_05408_),
    .A2(_05401_),
    .ZN(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11892_ (.I0(_05385_),
    .I1(\mod.u_cpu.rf_ram.memory[226][0] ),
    .S(_05409_),
    .Z(_05410_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11893_ (.I(_05410_),
    .Z(_00786_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11894_ (.I0(_05406_),
    .I1(\mod.u_cpu.rf_ram.memory[226][1] ),
    .S(_05409_),
    .Z(_05411_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11895_ (.I(_05411_),
    .Z(_00787_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11896_ (.I(_05309_),
    .Z(_05412_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11897_ (.I(_05412_),
    .Z(_05413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11898_ (.A1(_04973_),
    .A2(_05401_),
    .ZN(_05414_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11899_ (.I0(_05413_),
    .I1(\mod.u_cpu.rf_ram.memory[225][0] ),
    .S(_05414_),
    .Z(_05415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11900_ (.I(_05415_),
    .Z(_00788_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11901_ (.I0(_05406_),
    .I1(\mod.u_cpu.rf_ram.memory[225][1] ),
    .S(_05414_),
    .Z(_05416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11902_ (.I(_05416_),
    .Z(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11903_ (.I(_03984_),
    .Z(_05417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11904_ (.A1(_05417_),
    .A2(_05401_),
    .ZN(_05418_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11905_ (.I0(_05413_),
    .I1(\mod.u_cpu.rf_ram.memory[224][0] ),
    .S(_05418_),
    .Z(_05419_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11906_ (.I(_05419_),
    .Z(_00790_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11907_ (.I0(_05406_),
    .I1(\mod.u_cpu.rf_ram.memory[224][1] ),
    .S(_05418_),
    .Z(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11908_ (.I(_05420_),
    .Z(_00791_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11909_ (.A1(_04300_),
    .A2(_05371_),
    .ZN(_05421_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11910_ (.I(_05421_),
    .Z(_05422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11911_ (.I(_05422_),
    .Z(_05423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11912_ (.A1(_04845_),
    .A2(_05423_),
    .ZN(_05424_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11913_ (.I0(_05413_),
    .I1(\mod.u_cpu.rf_ram.memory[223][0] ),
    .S(_05424_),
    .Z(_05425_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11914_ (.I(_05425_),
    .Z(_00792_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11915_ (.I(_05405_),
    .Z(_05426_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11916_ (.I0(_05426_),
    .I1(\mod.u_cpu.rf_ram.memory[223][1] ),
    .S(_05424_),
    .Z(_05427_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11917_ (.I(_05427_),
    .Z(_00793_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11918_ (.I(_03750_),
    .Z(_05428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11919_ (.A1(_05428_),
    .A2(_05423_),
    .ZN(_05429_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11920_ (.I0(_05413_),
    .I1(\mod.u_cpu.rf_ram.memory[222][0] ),
    .S(_05429_),
    .Z(_05430_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11921_ (.I(_05430_),
    .Z(_00794_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11922_ (.I0(_05426_),
    .I1(\mod.u_cpu.rf_ram.memory[222][1] ),
    .S(_05429_),
    .Z(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11923_ (.I(_05431_),
    .Z(_00795_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11924_ (.I(_05421_),
    .Z(_05432_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11925_ (.I(_05432_),
    .Z(_05433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11926_ (.A1(_04994_),
    .A2(_05433_),
    .ZN(_05434_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11927_ (.A1(_05348_),
    .A2(_05434_),
    .ZN(_05435_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11928_ (.A1(_02192_),
    .A2(_05434_),
    .B(_05435_),
    .ZN(_00796_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11929_ (.I0(_05426_),
    .I1(\mod.u_cpu.rf_ram.memory[221][1] ),
    .S(_05434_),
    .Z(_05436_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11930_ (.I(_05436_),
    .Z(_00797_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11931_ (.I(_03698_),
    .Z(_05437_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11932_ (.A1(_03892_),
    .A2(_05319_),
    .ZN(_05438_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11933_ (.A1(_05078_),
    .A2(_05438_),
    .ZN(_05439_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11934_ (.I0(\mod.u_cpu.rf_ram.memory[169][0] ),
    .I1(_05437_),
    .S(_05439_),
    .Z(_05440_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11935_ (.I(_05440_),
    .Z(_00798_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11936_ (.I0(\mod.u_cpu.rf_ram.memory[169][1] ),
    .I1(_05230_),
    .S(_05439_),
    .Z(_05441_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11937_ (.I(_05441_),
    .Z(_00799_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11938_ (.I(_05412_),
    .Z(_05442_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11939_ (.I(_03780_),
    .Z(_05443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11940_ (.A1(_05443_),
    .A2(_05423_),
    .ZN(_05444_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11941_ (.I0(_05442_),
    .I1(\mod.u_cpu.rf_ram.memory[220][0] ),
    .S(_05444_),
    .Z(_05445_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11942_ (.I(_05445_),
    .Z(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11943_ (.I0(_05426_),
    .I1(\mod.u_cpu.rf_ram.memory[220][1] ),
    .S(_05444_),
    .Z(_05446_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11944_ (.I(_05446_),
    .Z(_00801_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11945_ (.A1(_04983_),
    .A2(_03837_),
    .ZN(_05447_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11946_ (.I(_05132_),
    .Z(_05448_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11947_ (.A1(_05448_),
    .A2(_05447_),
    .ZN(_05449_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11948_ (.A1(_02407_),
    .A2(_05447_),
    .B(_05449_),
    .ZN(_00802_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11949_ (.I(_05405_),
    .Z(_05450_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11950_ (.I0(_05450_),
    .I1(\mod.u_cpu.rf_ram.memory[21][1] ),
    .S(_05447_),
    .Z(_05451_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11951_ (.I(_05451_),
    .Z(_00803_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11952_ (.I(_03795_),
    .Z(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11953_ (.A1(_05452_),
    .A2(_05423_),
    .ZN(_05453_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11954_ (.I0(_05442_),
    .I1(\mod.u_cpu.rf_ram.memory[218][0] ),
    .S(_05453_),
    .Z(_05454_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11955_ (.I(_05454_),
    .Z(_00804_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11956_ (.I0(_05450_),
    .I1(\mod.u_cpu.rf_ram.memory[218][1] ),
    .S(_05453_),
    .Z(_05455_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11957_ (.I(_05455_),
    .Z(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11958_ (.A1(_05047_),
    .A2(_04118_),
    .ZN(_05456_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11959_ (.I0(_05442_),
    .I1(\mod.u_cpu.rf_ram.memory[529][0] ),
    .S(_05456_),
    .Z(_05457_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11960_ (.I(_05457_),
    .Z(_00806_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11961_ (.I0(_05450_),
    .I1(\mod.u_cpu.rf_ram.memory[529][1] ),
    .S(_05456_),
    .Z(_05458_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11962_ (.I(_05458_),
    .Z(_00807_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11963_ (.A1(_05139_),
    .A2(_03996_),
    .ZN(_05459_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11964_ (.I0(_05442_),
    .I1(\mod.u_cpu.rf_ram.memory[539][0] ),
    .S(_05459_),
    .Z(_05460_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11965_ (.I(_05460_),
    .Z(_00808_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11966_ (.I0(_05450_),
    .I1(\mod.u_cpu.rf_ram.memory[539][1] ),
    .S(_05459_),
    .Z(_05461_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11967_ (.I(_05461_),
    .Z(_00809_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11968_ (.A1(_04025_),
    .A2(_05433_),
    .ZN(_05462_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11969_ (.A1(_05448_),
    .A2(_05462_),
    .ZN(_05463_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11970_ (.A1(_02203_),
    .A2(_05462_),
    .B(_05463_),
    .ZN(_00810_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11971_ (.I(_05405_),
    .Z(_05464_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11972_ (.I0(_05464_),
    .I1(\mod.u_cpu.rf_ram.memory[217][1] ),
    .S(_05462_),
    .Z(_05465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11973_ (.I(_05465_),
    .Z(_00811_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11974_ (.A1(_03893_),
    .A2(_04108_),
    .ZN(_05466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11975_ (.A1(_05322_),
    .A2(_05466_),
    .ZN(_05467_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11976_ (.A1(_02458_),
    .A2(_05466_),
    .B(_05467_),
    .ZN(_00812_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11977_ (.I(_05229_),
    .Z(_05468_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11978_ (.I0(\mod.u_cpu.rf_ram.memory[549][1] ),
    .I1(_05468_),
    .S(_05466_),
    .Z(_05469_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11979_ (.I(_05469_),
    .Z(_00813_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11980_ (.I(_05412_),
    .Z(_05470_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11981_ (.I(_05422_),
    .Z(_05471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11982_ (.A1(_05283_),
    .A2(_05471_),
    .ZN(_05472_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11983_ (.I0(_05470_),
    .I1(\mod.u_cpu.rf_ram.memory[216][0] ),
    .S(_05472_),
    .Z(_05473_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11984_ (.I(_05473_),
    .Z(_00814_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11985_ (.I0(_05464_),
    .I1(\mod.u_cpu.rf_ram.memory[216][1] ),
    .S(_05472_),
    .Z(_05474_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11986_ (.I(_05474_),
    .Z(_00815_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11987_ (.A1(_03834_),
    .A2(_04068_),
    .ZN(_05475_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11988_ (.A1(_05448_),
    .A2(_05475_),
    .ZN(_05476_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11989_ (.A1(_02485_),
    .A2(_05475_),
    .B(_05476_),
    .ZN(_00816_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11990_ (.I0(_05464_),
    .I1(\mod.u_cpu.rf_ram.memory[559][1] ),
    .S(_05475_),
    .Z(_05477_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11991_ (.I(_05477_),
    .Z(_00817_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11992_ (.A1(_03767_),
    .A2(_04026_),
    .ZN(_05478_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11993_ (.I0(_05470_),
    .I1(\mod.u_cpu.rf_ram.memory[569][0] ),
    .S(_05478_),
    .Z(_05479_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11994_ (.I(_05479_),
    .Z(_00818_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11995_ (.I0(_05464_),
    .I1(\mod.u_cpu.rf_ram.memory[569][1] ),
    .S(_05478_),
    .Z(_05480_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11996_ (.I(_05480_),
    .Z(_00819_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11997_ (.A1(_05019_),
    .A2(_05433_),
    .ZN(_05481_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11998_ (.A1(_05448_),
    .A2(_05481_),
    .ZN(_05482_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11999_ (.A1(_02221_),
    .A2(_05481_),
    .B(_05482_),
    .ZN(_00820_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12000_ (.I(_05404_),
    .Z(_05483_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12001_ (.I(_05483_),
    .Z(_05484_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12002_ (.I0(_05484_),
    .I1(\mod.u_cpu.rf_ram.memory[215][1] ),
    .S(_05481_),
    .Z(_05485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12003_ (.I(_05485_),
    .Z(_00821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12004_ (.A1(_03834_),
    .A2(_04984_),
    .ZN(_05486_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12005_ (.I(_03773_),
    .Z(_05487_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12006_ (.I(_05487_),
    .Z(_05488_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12007_ (.A1(_05488_),
    .A2(_05486_),
    .ZN(_05489_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12008_ (.A1(_02501_),
    .A2(_05486_),
    .B(_05489_),
    .ZN(_00822_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12009_ (.I0(_05484_),
    .I1(\mod.u_cpu.rf_ram.memory[575][1] ),
    .S(_05486_),
    .Z(_05490_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12010_ (.I(_05490_),
    .Z(_00823_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12011_ (.A1(_04294_),
    .A2(_04026_),
    .ZN(_05491_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12012_ (.I0(_05470_),
    .I1(\mod.u_cpu.rf_ram.memory[57][0] ),
    .S(_05491_),
    .Z(_05492_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12013_ (.I(_05492_),
    .Z(_00824_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12014_ (.I0(_05484_),
    .I1(\mod.u_cpu.rf_ram.memory[57][1] ),
    .S(_05491_),
    .Z(_05493_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12015_ (.I(_05493_),
    .Z(_00825_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12016_ (.I(_03827_),
    .Z(_05494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12017_ (.A1(_05494_),
    .A2(_05471_),
    .ZN(_05495_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12018_ (.I0(_05470_),
    .I1(\mod.u_cpu.rf_ram.memory[214][0] ),
    .S(_05495_),
    .Z(_05496_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12019_ (.I(_05496_),
    .Z(_00826_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12020_ (.I0(_05484_),
    .I1(\mod.u_cpu.rf_ram.memory[214][1] ),
    .S(_05495_),
    .Z(_05497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12021_ (.I(_05497_),
    .Z(_00827_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12022_ (.I(_05412_),
    .Z(_05498_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12023_ (.A1(_05452_),
    .A2(_03810_),
    .ZN(_05499_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12024_ (.I0(_05498_),
    .I1(\mod.u_cpu.rf_ram.memory[58][0] ),
    .S(_05499_),
    .Z(_05500_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12025_ (.I(_05500_),
    .Z(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12026_ (.I(_05483_),
    .Z(_05501_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12027_ (.I0(_05501_),
    .I1(\mod.u_cpu.rf_ram.memory[58][1] ),
    .S(_05499_),
    .Z(_05502_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12028_ (.I(_05502_),
    .Z(_00829_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12029_ (.A1(_05239_),
    .A2(_03851_),
    .ZN(_05503_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12030_ (.I0(_05498_),
    .I1(\mod.u_cpu.rf_ram.memory[19][0] ),
    .S(_05503_),
    .Z(_05504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12031_ (.I(_05504_),
    .Z(_00830_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12032_ (.I0(_05501_),
    .I1(\mod.u_cpu.rf_ram.memory[19][1] ),
    .S(_05503_),
    .Z(_05505_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12033_ (.I(_05505_),
    .Z(_00831_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12034_ (.A1(_03728_),
    .A2(_04955_),
    .ZN(_05506_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12035_ (.I0(\mod.u_cpu.rf_ram.memory[5][0] ),
    .I1(_05437_),
    .S(_05506_),
    .Z(_05507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12036_ (.I(_05507_),
    .Z(_00832_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12037_ (.I0(\mod.u_cpu.rf_ram.memory[5][1] ),
    .I1(_05468_),
    .S(_05506_),
    .Z(_05508_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12038_ (.I(_05508_),
    .Z(_00833_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12039_ (.A1(_05443_),
    .A2(_03810_),
    .ZN(_05509_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12040_ (.I0(_05498_),
    .I1(\mod.u_cpu.rf_ram.memory[60][0] ),
    .S(_05509_),
    .Z(_05510_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12041_ (.I(_05510_),
    .Z(_00834_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12042_ (.I0(_05501_),
    .I1(\mod.u_cpu.rf_ram.memory[60][1] ),
    .S(_05509_),
    .Z(_05511_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12043_ (.I(_05511_),
    .Z(_00835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12044_ (.A1(_05164_),
    .A2(_05433_),
    .ZN(_05512_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12045_ (.A1(_05488_),
    .A2(_05512_),
    .ZN(_05513_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12046_ (.A1(_02226_),
    .A2(_05512_),
    .B(_05513_),
    .ZN(_00836_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12047_ (.I0(_05501_),
    .I1(\mod.u_cpu.rf_ram.memory[213][1] ),
    .S(_05512_),
    .Z(_05514_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12048_ (.I(_05514_),
    .Z(_00837_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12049_ (.I(_03770_),
    .Z(_05515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12050_ (.A1(_05515_),
    .A2(_03810_),
    .ZN(_05516_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12051_ (.I0(_05498_),
    .I1(\mod.u_cpu.rf_ram.memory[61][0] ),
    .S(_05516_),
    .Z(_05517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12052_ (.I(_05517_),
    .Z(_00838_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12053_ (.I(_05483_),
    .Z(_05518_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12054_ (.I0(_05518_),
    .I1(\mod.u_cpu.rf_ram.memory[61][1] ),
    .S(_05516_),
    .Z(_05519_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12055_ (.I(_05519_),
    .Z(_00839_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12056_ (.I(_05309_),
    .Z(_05520_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12057_ (.I(_05520_),
    .Z(_05521_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12058_ (.A1(_05428_),
    .A2(_03878_),
    .ZN(_05522_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12059_ (.I0(_05521_),
    .I1(\mod.u_cpu.rf_ram.memory[62][0] ),
    .S(_05522_),
    .Z(_05523_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12060_ (.I(_05523_),
    .Z(_00840_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12061_ (.I0(_05518_),
    .I1(\mod.u_cpu.rf_ram.memory[62][1] ),
    .S(_05522_),
    .Z(_05524_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12062_ (.I(_05524_),
    .Z(_00841_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12063_ (.A1(_04983_),
    .A2(_03771_),
    .ZN(_05525_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12064_ (.A1(_05488_),
    .A2(_05525_),
    .ZN(_05526_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12065_ (.A1(_02395_),
    .A2(_05525_),
    .B(_05526_),
    .ZN(_00842_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12066_ (.I0(_05518_),
    .I1(\mod.u_cpu.rf_ram.memory[29][1] ),
    .S(_05525_),
    .Z(_05527_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12067_ (.I(_05527_),
    .Z(_00843_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12068_ (.A1(_04294_),
    .A2(_04845_),
    .ZN(_05528_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12069_ (.I0(_05521_),
    .I1(\mod.u_cpu.rf_ram.memory[63][0] ),
    .S(_05528_),
    .Z(_05529_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12070_ (.I(_05529_),
    .Z(_00844_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12071_ (.I0(_05518_),
    .I1(\mod.u_cpu.rf_ram.memory[63][1] ),
    .S(_05528_),
    .Z(_05530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12072_ (.I(_05530_),
    .Z(_00845_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12073_ (.A1(_05417_),
    .A2(_05388_),
    .ZN(_05531_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12074_ (.I0(_05521_),
    .I1(\mod.u_cpu.rf_ram.memory[64][0] ),
    .S(_05531_),
    .Z(_05532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12075_ (.I(_05532_),
    .Z(_00846_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12076_ (.I(_05483_),
    .Z(_05533_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12077_ (.I0(_05533_),
    .I1(\mod.u_cpu.rf_ram.memory[64][1] ),
    .S(_05531_),
    .Z(_05534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12078_ (.I(_05534_),
    .Z(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12079_ (.I(_03841_),
    .Z(_05535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12080_ (.A1(_05535_),
    .A2(_05471_),
    .ZN(_05536_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12081_ (.I0(_05521_),
    .I1(\mod.u_cpu.rf_ram.memory[212][0] ),
    .S(_05536_),
    .Z(_05537_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12082_ (.I(_05537_),
    .Z(_00848_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12083_ (.I0(_05533_),
    .I1(\mod.u_cpu.rf_ram.memory[212][1] ),
    .S(_05536_),
    .Z(_05538_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12084_ (.I(_05538_),
    .Z(_00849_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12085_ (.I(_05520_),
    .Z(_05539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12086_ (.A1(_04973_),
    .A2(_05388_),
    .ZN(_05540_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12087_ (.I0(_05539_),
    .I1(\mod.u_cpu.rf_ram.memory[65][0] ),
    .S(_05540_),
    .Z(_05541_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12088_ (.I(_05541_),
    .Z(_00850_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12089_ (.I0(_05533_),
    .I1(\mod.u_cpu.rf_ram.memory[65][1] ),
    .S(_05540_),
    .Z(_05542_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12090_ (.I(_05542_),
    .Z(_00851_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12091_ (.I(_05387_),
    .Z(_05543_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12092_ (.A1(_05408_),
    .A2(_05543_),
    .ZN(_05544_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12093_ (.I0(_05539_),
    .I1(\mod.u_cpu.rf_ram.memory[66][0] ),
    .S(_05544_),
    .Z(_05545_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12094_ (.I(_05545_),
    .Z(_00852_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12095_ (.I0(_05533_),
    .I1(\mod.u_cpu.rf_ram.memory[66][1] ),
    .S(_05544_),
    .Z(_05546_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12096_ (.I(_05546_),
    .Z(_00853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12097_ (.A1(_04965_),
    .A2(_05543_),
    .ZN(_05547_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12098_ (.I0(_05539_),
    .I1(\mod.u_cpu.rf_ram.memory[67][0] ),
    .S(_05547_),
    .Z(_05548_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12099_ (.I(_05548_),
    .Z(_00854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12100_ (.I(_05404_),
    .Z(_05549_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12101_ (.I(_05549_),
    .Z(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12102_ (.I0(_05550_),
    .I1(\mod.u_cpu.rf_ram.memory[67][1] ),
    .S(_05547_),
    .Z(_05551_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12103_ (.I(_05551_),
    .Z(_00855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12104_ (.I(_05432_),
    .Z(_05552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12105_ (.A1(_03850_),
    .A2(_05552_),
    .ZN(_05553_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12106_ (.A1(_05488_),
    .A2(_05553_),
    .ZN(_05554_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12107_ (.A1(_02210_),
    .A2(_05553_),
    .B(_05554_),
    .ZN(_00856_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12108_ (.I0(_05550_),
    .I1(\mod.u_cpu.rf_ram.memory[211][1] ),
    .S(_05553_),
    .Z(_05555_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12109_ (.I(_05555_),
    .Z(_00857_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12110_ (.A1(_05367_),
    .A2(_05543_),
    .ZN(_05556_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12111_ (.I0(_05539_),
    .I1(\mod.u_cpu.rf_ram.memory[68][0] ),
    .S(_05556_),
    .Z(_05557_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12112_ (.I(_05557_),
    .Z(_00858_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12113_ (.I0(_05550_),
    .I1(\mod.u_cpu.rf_ram.memory[68][1] ),
    .S(_05556_),
    .Z(_05558_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12114_ (.I(_05558_),
    .Z(_00859_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12115_ (.I(_05520_),
    .Z(_05559_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12116_ (.A1(_05293_),
    .A2(_05471_),
    .ZN(_05560_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12117_ (.I0(_05559_),
    .I1(\mod.u_cpu.rf_ram.memory[210][0] ),
    .S(_05560_),
    .Z(_05561_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12118_ (.I(_05561_),
    .Z(_00860_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12119_ (.I0(_05550_),
    .I1(\mod.u_cpu.rf_ram.memory[210][1] ),
    .S(_05560_),
    .Z(_05562_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12120_ (.I(_05562_),
    .Z(_00861_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12121_ (.I(_04982_),
    .Z(_05563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12122_ (.A1(_05563_),
    .A2(_03843_),
    .ZN(_05564_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12123_ (.I0(_05559_),
    .I1(\mod.u_cpu.rf_ram.memory[20][0] ),
    .S(_05564_),
    .Z(_05565_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12124_ (.I(_05565_),
    .Z(_00862_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12125_ (.I(_05549_),
    .Z(_05566_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12126_ (.I0(_05566_),
    .I1(\mod.u_cpu.rf_ram.memory[20][1] ),
    .S(_05564_),
    .Z(_05567_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12127_ (.I(_05567_),
    .Z(_00863_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12128_ (.I(_05422_),
    .Z(_05568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12129_ (.A1(_05300_),
    .A2(_05568_),
    .ZN(_05569_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12130_ (.I0(_05559_),
    .I1(\mod.u_cpu.rf_ram.memory[208][0] ),
    .S(_05569_),
    .Z(_05570_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12131_ (.I(_05570_),
    .Z(_00864_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12132_ (.I0(_05566_),
    .I1(\mod.u_cpu.rf_ram.memory[208][1] ),
    .S(_05569_),
    .Z(_05571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12133_ (.I(_05571_),
    .Z(_00865_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12134_ (.A1(_05334_),
    .A2(_05543_),
    .ZN(_05572_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12135_ (.I0(_05559_),
    .I1(\mod.u_cpu.rf_ram.memory[74][0] ),
    .S(_05572_),
    .Z(_05573_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12136_ (.I(_05573_),
    .Z(_00866_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12137_ (.I0(_05566_),
    .I1(\mod.u_cpu.rf_ram.memory[74][1] ),
    .S(_05572_),
    .Z(_05574_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12138_ (.I(_05574_),
    .Z(_00867_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12139_ (.I(_05520_),
    .Z(_05575_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12140_ (.I(_05387_),
    .Z(_05576_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12141_ (.A1(_04930_),
    .A2(_05576_),
    .ZN(_05577_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12142_ (.I0(_05575_),
    .I1(\mod.u_cpu.rf_ram.memory[75][0] ),
    .S(_05577_),
    .Z(_05578_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12143_ (.I(_05578_),
    .Z(_00868_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12144_ (.I0(_05566_),
    .I1(\mod.u_cpu.rf_ram.memory[75][1] ),
    .S(_05577_),
    .Z(_05579_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12145_ (.I(_05579_),
    .Z(_00869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12146_ (.A1(_05187_),
    .A2(_05552_),
    .ZN(_05580_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12147_ (.I(_05487_),
    .Z(_05581_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12148_ (.A1(_05581_),
    .A2(_05580_),
    .ZN(_05582_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12149_ (.A1(_02181_),
    .A2(_05580_),
    .B(_05582_),
    .ZN(_00870_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12150_ (.I(_05549_),
    .Z(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12151_ (.I0(_05583_),
    .I1(\mod.u_cpu.rf_ram.memory[207][1] ),
    .S(_05580_),
    .Z(_05584_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12152_ (.I(_05584_),
    .Z(_00871_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12153_ (.A1(_05312_),
    .A2(_05568_),
    .ZN(_05585_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12154_ (.I0(_05575_),
    .I1(\mod.u_cpu.rf_ram.memory[206][0] ),
    .S(_05585_),
    .Z(_05586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12155_ (.I(_05586_),
    .Z(_00872_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12156_ (.I0(_05583_),
    .I1(\mod.u_cpu.rf_ram.memory[206][1] ),
    .S(_05585_),
    .Z(_05587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12157_ (.I(_05587_),
    .Z(_00873_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12158_ (.I(_03712_),
    .Z(_05588_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12159_ (.A1(_03727_),
    .A2(_04379_),
    .ZN(_05589_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12160_ (.A1(_05588_),
    .A2(_05589_),
    .ZN(_05590_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12161_ (.I0(\mod.u_cpu.rf_ram.memory[73][0] ),
    .I1(_05437_),
    .S(_05590_),
    .Z(_05591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12162_ (.I(_05591_),
    .Z(_00874_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12163_ (.I0(\mod.u_cpu.rf_ram.memory[73][1] ),
    .I1(_05468_),
    .S(_05590_),
    .Z(_05592_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12164_ (.I(_05592_),
    .Z(_00875_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12165_ (.I(_03894_),
    .Z(_05593_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12166_ (.A1(_04379_),
    .A2(_05319_),
    .ZN(_05594_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12167_ (.A1(_05593_),
    .A2(_05594_),
    .ZN(_05595_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12168_ (.A1(_05322_),
    .A2(_05595_),
    .ZN(_05596_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12169_ (.A1(_02176_),
    .A2(_05595_),
    .B(_05596_),
    .ZN(_00876_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12170_ (.I0(\mod.u_cpu.rf_ram.memory[205][1] ),
    .I1(_05468_),
    .S(_05595_),
    .Z(_05597_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12171_ (.I(_05597_),
    .Z(_00877_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12172_ (.A1(_05325_),
    .A2(_05576_),
    .ZN(_05598_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12173_ (.I0(_05575_),
    .I1(\mod.u_cpu.rf_ram.memory[76][0] ),
    .S(_05598_),
    .Z(_05599_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12174_ (.I(_05599_),
    .Z(_00878_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12175_ (.I0(_05583_),
    .I1(\mod.u_cpu.rf_ram.memory[76][1] ),
    .S(_05598_),
    .Z(_05600_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12176_ (.I(_05600_),
    .Z(_00879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12177_ (.A1(_05325_),
    .A2(_05568_),
    .ZN(_05601_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12178_ (.I0(_05575_),
    .I1(\mod.u_cpu.rf_ram.memory[204][0] ),
    .S(_05601_),
    .Z(_05602_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12179_ (.I(_05602_),
    .Z(_00880_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12180_ (.I0(_05583_),
    .I1(\mod.u_cpu.rf_ram.memory[204][1] ),
    .S(_05601_),
    .Z(_05603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12181_ (.I(_05603_),
    .Z(_00881_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12182_ (.I(_05309_),
    .Z(_05604_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12183_ (.I(_05604_),
    .Z(_05605_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12184_ (.I(_03909_),
    .Z(_05606_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12185_ (.A1(_05606_),
    .A2(_05568_),
    .ZN(_05607_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12186_ (.I0(_05605_),
    .I1(\mod.u_cpu.rf_ram.memory[203][0] ),
    .S(_05607_),
    .Z(_05608_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12187_ (.I(_05608_),
    .Z(_00882_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12188_ (.I(_05549_),
    .Z(_05609_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12189_ (.I0(_05609_),
    .I1(\mod.u_cpu.rf_ram.memory[203][1] ),
    .S(_05607_),
    .Z(_05610_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12190_ (.I(_05610_),
    .Z(_00883_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12191_ (.I(_05432_),
    .Z(_05611_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12192_ (.A1(_05334_),
    .A2(_05611_),
    .ZN(_05612_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12193_ (.I0(_05605_),
    .I1(\mod.u_cpu.rf_ram.memory[202][0] ),
    .S(_05612_),
    .Z(_05613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12194_ (.I(_05613_),
    .Z(_00884_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12195_ (.I0(_05609_),
    .I1(\mod.u_cpu.rf_ram.memory[202][1] ),
    .S(_05612_),
    .Z(_05614_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12196_ (.I(_05614_),
    .Z(_00885_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12197_ (.A1(_05588_),
    .A2(_05594_),
    .ZN(_05615_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12198_ (.I0(\mod.u_cpu.rf_ram.memory[201][0] ),
    .I1(_05437_),
    .S(_05615_),
    .Z(_05616_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12199_ (.I(_05616_),
    .Z(_00886_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12200_ (.I(_05229_),
    .Z(_05617_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12201_ (.I0(\mod.u_cpu.rf_ram.memory[201][1] ),
    .I1(_05617_),
    .S(_05615_),
    .Z(_05618_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12202_ (.I(_05618_),
    .Z(_00887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12203_ (.A1(_05343_),
    .A2(_05611_),
    .ZN(_05619_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12204_ (.I0(_05605_),
    .I1(\mod.u_cpu.rf_ram.memory[200][0] ),
    .S(_05619_),
    .Z(_05620_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12205_ (.I(_05620_),
    .Z(_00888_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12206_ (.I0(_05609_),
    .I1(\mod.u_cpu.rf_ram.memory[200][1] ),
    .S(_05619_),
    .Z(_05621_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12207_ (.I(_05621_),
    .Z(_00889_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12208_ (.I(_03698_),
    .Z(_05622_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12209_ (.A1(_04195_),
    .A2(_04125_),
    .Z(_05623_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12210_ (.I0(\mod.u_cpu.rf_ram.memory[1][0] ),
    .I1(_05622_),
    .S(_05623_),
    .Z(_05624_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12211_ (.I(_05624_),
    .Z(_00890_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12212_ (.I0(\mod.u_cpu.rf_ram.memory[1][1] ),
    .I1(_05617_),
    .S(_05623_),
    .Z(_05625_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12213_ (.I(_05625_),
    .Z(_00891_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12214_ (.A1(_05355_),
    .A2(_05611_),
    .ZN(_05626_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12215_ (.I0(_05605_),
    .I1(\mod.u_cpu.rf_ram.memory[198][0] ),
    .S(_05626_),
    .Z(_05627_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12216_ (.I(_05627_),
    .Z(_00892_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12217_ (.I0(_05609_),
    .I1(\mod.u_cpu.rf_ram.memory[198][1] ),
    .S(_05626_),
    .Z(_05628_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12218_ (.I(_05628_),
    .Z(_00893_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12219_ (.A1(_03726_),
    .A2(_04226_),
    .Z(_05629_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12220_ (.I(_05629_),
    .Z(_05630_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12221_ (.I(_05630_),
    .Z(_05631_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12222_ (.A1(_05019_),
    .A2(_05631_),
    .ZN(_05632_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12223_ (.A1(_05581_),
    .A2(_05632_),
    .ZN(_05633_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12224_ (.A1(_02330_),
    .A2(_05632_),
    .B(_05633_),
    .ZN(_00894_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12225_ (.I(_05404_),
    .Z(_05634_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12226_ (.I(_05634_),
    .Z(_05635_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12227_ (.I0(_05635_),
    .I1(\mod.u_cpu.rf_ram.memory[119][1] ),
    .S(_05632_),
    .Z(_05636_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12228_ (.I(_05636_),
    .Z(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12229_ (.A1(_05226_),
    .A2(_05594_),
    .ZN(_05637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12230_ (.A1(_05322_),
    .A2(_05637_),
    .ZN(_05638_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12231_ (.A1(_02158_),
    .A2(_05637_),
    .B(_05638_),
    .ZN(_00896_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12232_ (.I0(\mod.u_cpu.rf_ram.memory[197][1] ),
    .I1(_05617_),
    .S(_05637_),
    .Z(_05639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12233_ (.I(_05639_),
    .Z(_00897_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12234_ (.A1(_03727_),
    .A2(_04227_),
    .ZN(_05640_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12235_ (.A1(_05593_),
    .A2(_05640_),
    .ZN(_05641_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12236_ (.I(_03944_),
    .Z(_05642_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12237_ (.A1(_05642_),
    .A2(_05641_),
    .ZN(_05643_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12238_ (.A1(_02299_),
    .A2(_05641_),
    .B(_05643_),
    .ZN(_00898_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12239_ (.I0(\mod.u_cpu.rf_ram.memory[109][1] ),
    .I1(_05617_),
    .S(_05641_),
    .Z(_05644_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12240_ (.I(_05644_),
    .Z(_00899_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12241_ (.I(_05604_),
    .Z(_05645_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12242_ (.A1(_05367_),
    .A2(_05611_),
    .ZN(_05646_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12243_ (.I0(_05645_),
    .I1(\mod.u_cpu.rf_ram.memory[196][0] ),
    .S(_05646_),
    .Z(_05647_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12244_ (.I(_05647_),
    .Z(_00900_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12245_ (.I0(_05635_),
    .I1(\mod.u_cpu.rf_ram.memory[196][1] ),
    .S(_05646_),
    .Z(_05648_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12246_ (.I(_05648_),
    .Z(_00901_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _12247_ (.I(_03967_),
    .Z(_05649_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12248_ (.I(_05432_),
    .Z(_05650_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12249_ (.A1(_05649_),
    .A2(_05650_),
    .ZN(_05651_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12250_ (.I0(_05645_),
    .I1(\mod.u_cpu.rf_ram.memory[195][0] ),
    .S(_05651_),
    .Z(_05652_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12251_ (.I(_05652_),
    .Z(_00902_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12252_ (.I0(_05635_),
    .I1(\mod.u_cpu.rf_ram.memory[195][1] ),
    .S(_05651_),
    .Z(_05653_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12253_ (.I(_05653_),
    .Z(_00903_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12254_ (.A1(_05408_),
    .A2(_05650_),
    .ZN(_05654_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12255_ (.I0(_05645_),
    .I1(\mod.u_cpu.rf_ram.memory[194][0] ),
    .S(_05654_),
    .Z(_05655_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12256_ (.I(_05655_),
    .Z(_00904_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12257_ (.I0(_05635_),
    .I1(\mod.u_cpu.rf_ram.memory[194][1] ),
    .S(_05654_),
    .Z(_05656_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12258_ (.I(_05656_),
    .Z(_00905_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12259_ (.I(_03979_),
    .Z(_05657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12260_ (.A1(_05657_),
    .A2(_05650_),
    .ZN(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12261_ (.I0(_05645_),
    .I1(\mod.u_cpu.rf_ram.memory[193][0] ),
    .S(_05658_),
    .Z(_05659_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12262_ (.I(_05659_),
    .Z(_00906_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12263_ (.I(_05634_),
    .Z(_05660_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12264_ (.I0(_05660_),
    .I1(\mod.u_cpu.rf_ram.memory[193][1] ),
    .S(_05658_),
    .Z(_05661_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12265_ (.I(_05661_),
    .Z(_00907_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12266_ (.I(_05604_),
    .Z(_05662_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12267_ (.A1(_05417_),
    .A2(_05650_),
    .ZN(_05663_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12268_ (.I0(_05662_),
    .I1(\mod.u_cpu.rf_ram.memory[192][0] ),
    .S(_05663_),
    .Z(_05664_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12269_ (.I(_05664_),
    .Z(_00908_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12270_ (.I0(_05660_),
    .I1(\mod.u_cpu.rf_ram.memory[192][1] ),
    .S(_05663_),
    .Z(_05665_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12271_ (.I(_05665_),
    .Z(_00909_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12272_ (.A1(_03755_),
    .A2(_05371_),
    .ZN(_05666_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12273_ (.I(_05666_),
    .Z(_05667_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12274_ (.I(_05667_),
    .Z(_05668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12275_ (.A1(_04984_),
    .A2(_05668_),
    .ZN(_05669_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12276_ (.I0(_05662_),
    .I1(\mod.u_cpu.rf_ram.memory[191][0] ),
    .S(_05669_),
    .Z(_05670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12277_ (.I(_05670_),
    .Z(_00910_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12278_ (.I0(_05660_),
    .I1(\mod.u_cpu.rf_ram.memory[191][1] ),
    .S(_05669_),
    .Z(_05671_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12279_ (.I(_05671_),
    .Z(_00911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12280_ (.A1(_05428_),
    .A2(_05668_),
    .ZN(_05672_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12281_ (.I0(_05662_),
    .I1(\mod.u_cpu.rf_ram.memory[190][0] ),
    .S(_05672_),
    .Z(_05673_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12282_ (.I(_05673_),
    .Z(_00912_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12283_ (.I0(_05660_),
    .I1(\mod.u_cpu.rf_ram.memory[190][1] ),
    .S(_05672_),
    .Z(_05674_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12284_ (.I(_05674_),
    .Z(_00913_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12285_ (.A1(_05563_),
    .A2(_03859_),
    .ZN(_05675_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12286_ (.I0(_05662_),
    .I1(\mod.u_cpu.rf_ram.memory[18][0] ),
    .S(_05675_),
    .Z(_05676_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12287_ (.I(_05676_),
    .Z(_00914_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12288_ (.I(_05634_),
    .Z(_05677_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12289_ (.I0(_05677_),
    .I1(\mod.u_cpu.rf_ram.memory[18][1] ),
    .S(_05675_),
    .Z(_05678_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12290_ (.I(_05678_),
    .Z(_00915_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12291_ (.I(_05604_),
    .Z(_05679_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12292_ (.A1(_05443_),
    .A2(_05668_),
    .ZN(_05680_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12293_ (.I0(_05679_),
    .I1(\mod.u_cpu.rf_ram.memory[188][0] ),
    .S(_05680_),
    .Z(_05681_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12294_ (.I(_05681_),
    .Z(_00916_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12295_ (.I0(_05677_),
    .I1(\mod.u_cpu.rf_ram.memory[188][1] ),
    .S(_05680_),
    .Z(_05682_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12296_ (.I(_05682_),
    .Z(_00917_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12297_ (.A1(_05139_),
    .A2(_05668_),
    .ZN(_05683_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12298_ (.I0(_05679_),
    .I1(\mod.u_cpu.rf_ram.memory[187][0] ),
    .S(_05683_),
    .Z(_05684_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12299_ (.I(_05684_),
    .Z(_00918_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12300_ (.I0(_05677_),
    .I1(\mod.u_cpu.rf_ram.memory[187][1] ),
    .S(_05683_),
    .Z(_05685_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12301_ (.I(_05685_),
    .Z(_00919_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12302_ (.I(_05667_),
    .Z(_05686_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12303_ (.A1(_05452_),
    .A2(_05686_),
    .ZN(_05687_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12304_ (.I0(_05679_),
    .I1(\mod.u_cpu.rf_ram.memory[186][0] ),
    .S(_05687_),
    .Z(_05688_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12305_ (.I(_05688_),
    .Z(_00920_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12306_ (.I0(_05677_),
    .I1(\mod.u_cpu.rf_ram.memory[186][1] ),
    .S(_05687_),
    .Z(_05689_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12307_ (.I(_05689_),
    .Z(_00921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12308_ (.A1(_04873_),
    .A2(_05686_),
    .ZN(_05690_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12309_ (.I0(_05679_),
    .I1(\mod.u_cpu.rf_ram.memory[185][0] ),
    .S(_05690_),
    .Z(_05691_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12310_ (.I(_05691_),
    .Z(_00922_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12311_ (.I(_05634_),
    .Z(_05692_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12312_ (.I0(_05692_),
    .I1(\mod.u_cpu.rf_ram.memory[185][1] ),
    .S(_05690_),
    .Z(_05693_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12313_ (.I(_05693_),
    .Z(_00923_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12314_ (.I(_03696_),
    .Z(_05694_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12315_ (.I(_05694_),
    .Z(_05695_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12316_ (.I(_05695_),
    .Z(_05696_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12317_ (.A1(_05515_),
    .A2(_05686_),
    .ZN(_05697_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12318_ (.I0(_05696_),
    .I1(\mod.u_cpu.rf_ram.memory[189][0] ),
    .S(_05697_),
    .Z(_05698_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12319_ (.I(_05698_),
    .Z(_00924_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12320_ (.I0(_05692_),
    .I1(\mod.u_cpu.rf_ram.memory[189][1] ),
    .S(_05697_),
    .Z(_05699_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12321_ (.I(_05699_),
    .Z(_00925_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12322_ (.A1(_05037_),
    .A2(_05686_),
    .ZN(_05700_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12323_ (.I0(_05696_),
    .I1(\mod.u_cpu.rf_ram.memory[179][0] ),
    .S(_05700_),
    .Z(_05701_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12324_ (.I(_05701_),
    .Z(_00926_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12325_ (.I0(_05692_),
    .I1(\mod.u_cpu.rf_ram.memory[179][1] ),
    .S(_05700_),
    .Z(_05702_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12326_ (.I(_05702_),
    .Z(_00927_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12327_ (.I(_05667_),
    .Z(_05703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12328_ (.A1(_05283_),
    .A2(_05703_),
    .ZN(_05704_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12329_ (.I0(_05696_),
    .I1(\mod.u_cpu.rf_ram.memory[184][0] ),
    .S(_05704_),
    .Z(_05705_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12330_ (.I(_05705_),
    .Z(_00928_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12331_ (.I0(_05692_),
    .I1(\mod.u_cpu.rf_ram.memory[184][1] ),
    .S(_05704_),
    .Z(_05706_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12332_ (.I(_05706_),
    .Z(_00929_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12333_ (.A1(_03879_),
    .A2(_05703_),
    .ZN(_05707_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12334_ (.I0(_05696_),
    .I1(\mod.u_cpu.rf_ram.memory[183][0] ),
    .S(_05707_),
    .Z(_05708_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12335_ (.I(_05708_),
    .Z(_00930_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12336_ (.I(_05105_),
    .Z(_05709_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12337_ (.I(_05709_),
    .Z(_05710_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12338_ (.I(_05710_),
    .Z(_05711_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12339_ (.I0(_05711_),
    .I1(\mod.u_cpu.rf_ram.memory[183][1] ),
    .S(_05707_),
    .Z(_05712_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12340_ (.I(_05712_),
    .Z(_00931_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12341_ (.I(_05695_),
    .Z(_05713_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12342_ (.A1(_05494_),
    .A2(_05703_),
    .ZN(_05714_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12343_ (.I0(_05713_),
    .I1(\mod.u_cpu.rf_ram.memory[182][0] ),
    .S(_05714_),
    .Z(_05715_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12344_ (.I(_05715_),
    .Z(_00932_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12345_ (.I0(_05711_),
    .I1(\mod.u_cpu.rf_ram.memory[182][1] ),
    .S(_05714_),
    .Z(_05716_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12346_ (.I(_05716_),
    .Z(_00933_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12347_ (.A1(_04014_),
    .A2(_05703_),
    .ZN(_05717_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12348_ (.I0(_05713_),
    .I1(\mod.u_cpu.rf_ram.memory[181][0] ),
    .S(_05717_),
    .Z(_05718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12349_ (.I(_05718_),
    .Z(_00934_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12350_ (.I0(_05711_),
    .I1(\mod.u_cpu.rf_ram.memory[181][1] ),
    .S(_05717_),
    .Z(_05719_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12351_ (.I(_05719_),
    .Z(_00935_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12352_ (.I(_05629_),
    .Z(_05720_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12353_ (.I(_05720_),
    .Z(_05721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12354_ (.A1(_05452_),
    .A2(_05721_),
    .ZN(_05722_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12355_ (.I0(_05713_),
    .I1(\mod.u_cpu.rf_ram.memory[122][0] ),
    .S(_05722_),
    .Z(_05723_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12356_ (.I(_05723_),
    .Z(_00936_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12357_ (.I0(_05711_),
    .I1(\mod.u_cpu.rf_ram.memory[122][1] ),
    .S(_05722_),
    .Z(_05724_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12358_ (.I(_05724_),
    .Z(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12359_ (.I(_05666_),
    .Z(_05725_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12360_ (.I(_05725_),
    .Z(_05726_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12361_ (.A1(_05535_),
    .A2(_05726_),
    .ZN(_05727_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12362_ (.I0(_05713_),
    .I1(\mod.u_cpu.rf_ram.memory[180][0] ),
    .S(_05727_),
    .Z(_05728_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12363_ (.I(_05728_),
    .Z(_00938_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12364_ (.I(_05710_),
    .Z(_05729_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12365_ (.I0(_05729_),
    .I1(\mod.u_cpu.rf_ram.memory[180][1] ),
    .S(_05727_),
    .Z(_05730_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12366_ (.I(_05730_),
    .Z(_00939_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12367_ (.I(_05695_),
    .Z(_05731_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12368_ (.I(_03849_),
    .Z(_05732_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12369_ (.A1(_05732_),
    .A2(_04137_),
    .ZN(_05733_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12370_ (.I0(_05731_),
    .I1(\mod.u_cpu.rf_ram.memory[499][0] ),
    .S(_05733_),
    .Z(_05734_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12371_ (.I(_05734_),
    .Z(_00940_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12372_ (.I0(_05729_),
    .I1(\mod.u_cpu.rf_ram.memory[499][1] ),
    .S(_05733_),
    .Z(_05735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12373_ (.I(_05735_),
    .Z(_00941_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12374_ (.A1(_05563_),
    .A2(_03866_),
    .ZN(_05736_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12375_ (.I0(_05731_),
    .I1(\mod.u_cpu.rf_ram.memory[17][0] ),
    .S(_05736_),
    .Z(_05737_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12376_ (.I(_05737_),
    .Z(_00942_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12377_ (.I0(_05729_),
    .I1(\mod.u_cpu.rf_ram.memory[17][1] ),
    .S(_05736_),
    .Z(_05738_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12378_ (.I(_05738_),
    .Z(_00943_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12379_ (.A1(_05293_),
    .A2(_05726_),
    .ZN(_05739_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12380_ (.I0(_05731_),
    .I1(\mod.u_cpu.rf_ram.memory[178][0] ),
    .S(_05739_),
    .Z(_05740_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12381_ (.I(_05740_),
    .Z(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12382_ (.I0(_05729_),
    .I1(\mod.u_cpu.rf_ram.memory[178][1] ),
    .S(_05739_),
    .Z(_05741_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12383_ (.I(_05741_),
    .Z(_00945_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12384_ (.I(_03864_),
    .Z(_05742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12385_ (.A1(_05742_),
    .A2(_05726_),
    .ZN(_05743_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12386_ (.I0(_05731_),
    .I1(\mod.u_cpu.rf_ram.memory[177][0] ),
    .S(_05743_),
    .Z(_05744_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12387_ (.I(_05744_),
    .Z(_00946_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12388_ (.I(_05710_),
    .Z(_05745_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12389_ (.I0(_05745_),
    .I1(\mod.u_cpu.rf_ram.memory[177][1] ),
    .S(_05743_),
    .Z(_05746_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12390_ (.I(_05746_),
    .Z(_00947_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12391_ (.A1(_03770_),
    .A2(_04142_),
    .ZN(_05747_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12392_ (.A1(_05581_),
    .A2(_05747_),
    .ZN(_05748_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12393_ (.A1(_01609_),
    .A2(_05747_),
    .B(_05748_),
    .ZN(_00948_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12394_ (.I0(_05745_),
    .I1(\mod.u_cpu.rf_ram.memory[509][1] ),
    .S(_05747_),
    .Z(_05749_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12395_ (.I(_05749_),
    .Z(_00949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12396_ (.A1(_04700_),
    .A2(_04335_),
    .ZN(_05750_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12397_ (.A1(_05581_),
    .A2(_05750_),
    .ZN(_05751_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12398_ (.A1(_01562_),
    .A2(_05750_),
    .B(_05751_),
    .ZN(_00950_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12399_ (.I0(_05745_),
    .I1(\mod.u_cpu.rf_ram.memory[479][1] ),
    .S(_05750_),
    .Z(_05752_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12400_ (.I(_05752_),
    .Z(_00951_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12401_ (.I(_05695_),
    .Z(_05753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12402_ (.A1(_05300_),
    .A2(_05726_),
    .ZN(_05754_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12403_ (.I0(_05753_),
    .I1(\mod.u_cpu.rf_ram.memory[176][0] ),
    .S(_05754_),
    .Z(_05755_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12404_ (.I(_05755_),
    .Z(_00952_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12405_ (.I0(_05745_),
    .I1(\mod.u_cpu.rf_ram.memory[176][1] ),
    .S(_05754_),
    .Z(_05756_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12406_ (.I(_05756_),
    .Z(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12407_ (.I(_05725_),
    .Z(_05757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12408_ (.A1(_05187_),
    .A2(_05757_),
    .ZN(_05758_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12409_ (.I(_05487_),
    .Z(_05759_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12410_ (.A1(_05759_),
    .A2(_05758_),
    .ZN(_05760_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12411_ (.A1(_02117_),
    .A2(_05758_),
    .B(_05760_),
    .ZN(_00954_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12412_ (.I(_05710_),
    .Z(_05761_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12413_ (.I0(_05761_),
    .I1(\mod.u_cpu.rf_ram.memory[175][1] ),
    .S(_05758_),
    .Z(_05762_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12414_ (.I(_05762_),
    .Z(_00955_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12415_ (.A1(_05588_),
    .A2(_04228_),
    .ZN(_05763_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12416_ (.I0(\mod.u_cpu.rf_ram.memory[489][0] ),
    .I1(_05622_),
    .S(_05763_),
    .Z(_05764_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12417_ (.I(_05764_),
    .Z(_00956_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12418_ (.I(_05229_),
    .Z(_05765_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12419_ (.I0(\mod.u_cpu.rf_ram.memory[489][1] ),
    .I1(_05765_),
    .S(_05763_),
    .Z(_05766_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12420_ (.I(_05766_),
    .Z(_00957_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12421_ (.I(_05725_),
    .Z(_05767_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12422_ (.A1(_05312_),
    .A2(_05767_),
    .ZN(_05768_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12423_ (.I0(_05753_),
    .I1(\mod.u_cpu.rf_ram.memory[174][0] ),
    .S(_05768_),
    .Z(_05769_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12424_ (.I(_05769_),
    .Z(_00958_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12425_ (.I0(_05761_),
    .I1(\mod.u_cpu.rf_ram.memory[174][1] ),
    .S(_05768_),
    .Z(_05770_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12426_ (.I(_05770_),
    .Z(_00959_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12427_ (.A1(_05019_),
    .A2(_04442_),
    .ZN(_05771_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12428_ (.A1(_05759_),
    .A2(_05771_),
    .ZN(_05772_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12429_ (.A1(_01796_),
    .A2(_05771_),
    .B(_05772_),
    .ZN(_00960_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12430_ (.I0(_05761_),
    .I1(\mod.u_cpu.rf_ram.memory[439][1] ),
    .S(_05771_),
    .Z(_05773_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12431_ (.I(_05773_),
    .Z(_00961_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12432_ (.A1(_05593_),
    .A2(_05438_),
    .ZN(_05774_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12433_ (.A1(_05642_),
    .A2(_05774_),
    .ZN(_05775_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12434_ (.A1(_02112_),
    .A2(_05774_),
    .B(_05775_),
    .ZN(_00962_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12435_ (.I0(\mod.u_cpu.rf_ram.memory[173][1] ),
    .I1(_05765_),
    .S(_05774_),
    .Z(_05776_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12436_ (.I(_05776_),
    .Z(_00963_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12437_ (.A1(_05325_),
    .A2(_05767_),
    .ZN(_05777_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12438_ (.I0(_05753_),
    .I1(\mod.u_cpu.rf_ram.memory[172][0] ),
    .S(_05777_),
    .Z(_05778_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12439_ (.I(_05778_),
    .Z(_00964_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12440_ (.I0(_05761_),
    .I1(\mod.u_cpu.rf_ram.memory[172][1] ),
    .S(_05777_),
    .Z(_05779_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12441_ (.I(_05779_),
    .Z(_00965_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12442_ (.I(_01433_),
    .Z(_05780_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12443_ (.I(_03498_),
    .Z(_05781_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _12444_ (.I(_05781_),
    .ZN(_05782_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12445_ (.I(_05782_),
    .Z(_05783_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12446_ (.I(_05783_),
    .Z(_05784_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12447_ (.A1(_03412_),
    .A2(_03400_),
    .ZN(_05785_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12448_ (.A1(\mod.u_arbiter.i_wb_cpu_ibus_adr[1] ),
    .A2(_05784_),
    .B(_05785_),
    .ZN(_05786_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12449_ (.I(_05786_),
    .Z(_05787_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12450_ (.A1(_05780_),
    .A2(\mod.u_cpu.cpu.state.stage_two_req ),
    .B(_05787_),
    .ZN(_05788_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12451_ (.A1(_03700_),
    .A2(_05788_),
    .ZN(_05789_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12452_ (.I(_03394_),
    .Z(_05790_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12453_ (.A1(_03289_),
    .A2(_03667_),
    .Z(_05791_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12454_ (.A1(_03281_),
    .A2(_05791_),
    .ZN(_05792_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _12455_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[2] ),
    .A2(_03430_),
    .A3(\mod.u_arbiter.i_wb_cpu_dbus_dat[1] ),
    .Z(_05793_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _12456_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[3] ),
    .A2(_05793_),
    .Z(_05794_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12457_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[4] ),
    .A2(_05794_),
    .ZN(_05795_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12458_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .A2(_05795_),
    .Z(_05796_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _12459_ (.A1(_03338_),
    .A2(_03668_),
    .B(_03359_),
    .C(_03394_),
    .ZN(_05797_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _12460_ (.A1(_05792_),
    .A2(_05796_),
    .B1(_05797_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[6] ),
    .ZN(_05798_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12461_ (.A1(_03359_),
    .A2(_03355_),
    .A3(_05798_),
    .ZN(_05799_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12462_ (.A1(\mod.u_arbiter.i_wb_cpu_ack ),
    .A2(_03406_),
    .Z(_05800_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12463_ (.I(_05800_),
    .Z(_05801_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _12464_ (.A1(_05790_),
    .A2(_05799_),
    .B(_05801_),
    .C(_03686_),
    .ZN(_05802_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _12465_ (.A1(_01433_),
    .A2(_03284_),
    .A3(_03377_),
    .A4(_05802_),
    .Z(_05803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12466_ (.A1(_05789_),
    .A2(_05803_),
    .ZN(_00966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12467_ (.A1(_05649_),
    .A2(_04437_),
    .ZN(_05804_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12468_ (.I0(_05753_),
    .I1(\mod.u_cpu.rf_ram.memory[419][0] ),
    .S(_05804_),
    .Z(_05805_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12469_ (.I(_05805_),
    .Z(_00967_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12470_ (.I(_05709_),
    .Z(_05806_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12471_ (.I(_05806_),
    .Z(_05807_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12472_ (.I0(_05807_),
    .I1(\mod.u_cpu.rf_ram.memory[419][1] ),
    .S(_05804_),
    .Z(_05808_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12473_ (.I(_05808_),
    .Z(_00968_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12474_ (.A1(_05395_),
    .A2(_04033_),
    .ZN(_05809_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12475_ (.A1(_05759_),
    .A2(_05809_),
    .ZN(_05810_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12476_ (.A1(_02535_),
    .A2(_05809_),
    .B(_05810_),
    .ZN(_00969_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12477_ (.I0(_05807_),
    .I1(\mod.u_cpu.rf_ram.memory[519][1] ),
    .S(_05809_),
    .Z(_05811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12478_ (.I(_05811_),
    .Z(_00970_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12479_ (.I(_05694_),
    .Z(_05812_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12480_ (.I(_05812_),
    .Z(_05813_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12481_ (.A1(_05657_),
    .A2(_04309_),
    .ZN(_05814_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12482_ (.I0(_05813_),
    .I1(\mod.u_cpu.rf_ram.memory[449][0] ),
    .S(_05814_),
    .Z(_05815_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12483_ (.I(_05815_),
    .Z(_00971_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12484_ (.I0(_05807_),
    .I1(\mod.u_cpu.rf_ram.memory[449][1] ),
    .S(_05814_),
    .Z(_05816_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12485_ (.I(_05816_),
    .Z(_00972_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12486_ (.A1(_05606_),
    .A2(_05767_),
    .ZN(_05817_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12487_ (.I0(_05813_),
    .I1(\mod.u_cpu.rf_ram.memory[171][0] ),
    .S(_05817_),
    .Z(_05818_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12488_ (.I(_05818_),
    .Z(_00973_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12489_ (.I0(_05807_),
    .I1(\mod.u_cpu.rf_ram.memory[171][1] ),
    .S(_05817_),
    .Z(_05819_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12490_ (.I(_05819_),
    .Z(_00974_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12491_ (.A1(_05334_),
    .A2(_05767_),
    .ZN(_05820_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12492_ (.I0(_05813_),
    .I1(\mod.u_cpu.rf_ram.memory[170][0] ),
    .S(_05820_),
    .Z(_05821_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12493_ (.I(_05821_),
    .Z(_00975_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12494_ (.I(_05806_),
    .Z(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12495_ (.I0(_05822_),
    .I1(\mod.u_cpu.rf_ram.memory[170][1] ),
    .S(_05820_),
    .Z(_05823_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12496_ (.I(_05823_),
    .Z(_00976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12497_ (.A1(_05606_),
    .A2(_04309_),
    .ZN(_05824_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12498_ (.I0(_05813_),
    .I1(\mod.u_cpu.rf_ram.memory[459][0] ),
    .S(_05824_),
    .Z(_05825_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12499_ (.I(_05825_),
    .Z(_00977_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12500_ (.I0(_05822_),
    .I1(\mod.u_cpu.rf_ram.memory[459][1] ),
    .S(_05824_),
    .Z(_05826_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12501_ (.I(_05826_),
    .Z(_00978_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12502_ (.I(_05812_),
    .Z(_05827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12503_ (.A1(_05563_),
    .A2(_03873_),
    .ZN(_05828_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12504_ (.I0(_05827_),
    .I1(\mod.u_cpu.rf_ram.memory[16][0] ),
    .S(_05828_),
    .Z(_05829_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12505_ (.I(_05829_),
    .Z(_00979_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12506_ (.I0(_05822_),
    .I1(\mod.u_cpu.rf_ram.memory[16][1] ),
    .S(_05828_),
    .Z(_05830_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12507_ (.I(_05830_),
    .Z(_00980_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12508_ (.I(_05725_),
    .Z(_05831_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12509_ (.A1(_05343_),
    .A2(_05831_),
    .ZN(_05832_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12510_ (.I0(_05827_),
    .I1(\mod.u_cpu.rf_ram.memory[168][0] ),
    .S(_05832_),
    .Z(_05833_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12511_ (.I(_05833_),
    .Z(_00981_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12512_ (.I0(_05822_),
    .I1(\mod.u_cpu.rf_ram.memory[168][1] ),
    .S(_05832_),
    .Z(_05834_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12513_ (.I(_05834_),
    .Z(_00982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12514_ (.A1(_05395_),
    .A2(_05667_),
    .ZN(_05835_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12515_ (.A1(_05759_),
    .A2(_05835_),
    .ZN(_05836_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12516_ (.A1(_02137_),
    .A2(_05835_),
    .B(_05836_),
    .ZN(_00983_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12517_ (.I(_05806_),
    .Z(_05837_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12518_ (.I0(_05837_),
    .I1(\mod.u_cpu.rf_ram.memory[167][1] ),
    .S(_05835_),
    .Z(_05838_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12519_ (.I(_05838_),
    .Z(_00984_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12520_ (.A1(_05355_),
    .A2(_05831_),
    .ZN(_05839_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12521_ (.I0(_05827_),
    .I1(\mod.u_cpu.rf_ram.memory[166][0] ),
    .S(_05839_),
    .Z(_05840_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12522_ (.I(_05840_),
    .Z(_00985_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12523_ (.I0(_05837_),
    .I1(\mod.u_cpu.rf_ram.memory[166][1] ),
    .S(_05839_),
    .Z(_05841_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12524_ (.I(_05841_),
    .Z(_00986_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12525_ (.A1(_05164_),
    .A2(_04302_),
    .ZN(_05842_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12526_ (.I(_05487_),
    .Z(_05843_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12527_ (.A1(_05843_),
    .A2(_05842_),
    .ZN(_05844_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12528_ (.A1(_01574_),
    .A2(_05842_),
    .B(_05844_),
    .ZN(_00987_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12529_ (.I0(_05837_),
    .I1(\mod.u_cpu.rf_ram.memory[469][1] ),
    .S(_05842_),
    .Z(_05845_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12530_ (.I(_05845_),
    .Z(_00988_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12531_ (.A1(_05593_),
    .A2(_04528_),
    .ZN(_05846_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12532_ (.A1(_05642_),
    .A2(_05846_),
    .ZN(_05847_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12533_ (.A1(_01775_),
    .A2(_05846_),
    .B(_05847_),
    .ZN(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12534_ (.I0(\mod.u_cpu.rf_ram.memory[429][1] ),
    .I1(_05765_),
    .S(_05846_),
    .Z(_05848_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12535_ (.I(_05848_),
    .Z(_00990_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12536_ (.A1(_05226_),
    .A2(_05438_),
    .ZN(_05849_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12537_ (.A1(_05642_),
    .A2(_05849_),
    .ZN(_05850_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12538_ (.A1(_02131_),
    .A2(_05849_),
    .B(_05850_),
    .ZN(_00991_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12539_ (.I0(\mod.u_cpu.rf_ram.memory[165][1] ),
    .I1(_05765_),
    .S(_05849_),
    .Z(_05851_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12540_ (.I(_05851_),
    .Z(_00992_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12541_ (.A1(_05367_),
    .A2(_05831_),
    .ZN(_05852_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12542_ (.I0(_05827_),
    .I1(\mod.u_cpu.rf_ram.memory[164][0] ),
    .S(_05852_),
    .Z(_05853_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12543_ (.I(_05853_),
    .Z(_00993_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12544_ (.I0(_05837_),
    .I1(\mod.u_cpu.rf_ram.memory[164][1] ),
    .S(_05852_),
    .Z(_05854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12545_ (.I(_05854_),
    .Z(_00994_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12546_ (.I(_05812_),
    .Z(_05855_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12547_ (.A1(_05649_),
    .A2(_05831_),
    .ZN(_05856_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12548_ (.I0(_05855_),
    .I1(\mod.u_cpu.rf_ram.memory[163][0] ),
    .S(_05856_),
    .Z(_05857_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12549_ (.I(_05857_),
    .Z(_00995_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12550_ (.I(_05806_),
    .Z(_05858_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12551_ (.I0(_05858_),
    .I1(\mod.u_cpu.rf_ram.memory[163][1] ),
    .S(_05856_),
    .Z(_05859_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12552_ (.I(_05859_),
    .Z(_00996_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12553_ (.A1(_05408_),
    .A2(_05757_),
    .ZN(_05860_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12554_ (.I0(_05855_),
    .I1(\mod.u_cpu.rf_ram.memory[162][0] ),
    .S(_05860_),
    .Z(_05861_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12555_ (.I(_05861_),
    .Z(_00997_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12556_ (.I0(_05858_),
    .I1(\mod.u_cpu.rf_ram.memory[162][1] ),
    .S(_05860_),
    .Z(_05862_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12557_ (.I(_05862_),
    .Z(_00998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12558_ (.A1(_05657_),
    .A2(_05757_),
    .ZN(_05863_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12559_ (.I0(_05855_),
    .I1(\mod.u_cpu.rf_ram.memory[161][0] ),
    .S(_05863_),
    .Z(_05864_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12560_ (.I(_05864_),
    .Z(_00999_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12561_ (.I0(_05858_),
    .I1(\mod.u_cpu.rf_ram.memory[161][1] ),
    .S(_05863_),
    .Z(_05865_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12562_ (.I(_05865_),
    .Z(_01000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12563_ (.A1(_05417_),
    .A2(_05757_),
    .ZN(_05866_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12564_ (.I0(_05855_),
    .I1(\mod.u_cpu.rf_ram.memory[160][0] ),
    .S(_05866_),
    .Z(_05867_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12565_ (.I(_05867_),
    .Z(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12566_ (.I0(_05858_),
    .I1(\mod.u_cpu.rf_ram.memory[160][1] ),
    .S(_05866_),
    .Z(_05868_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12567_ (.I(_05868_),
    .Z(_01002_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12568_ (.I(_05812_),
    .Z(_05869_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12569_ (.I(_04982_),
    .Z(_05870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12570_ (.A1(_05870_),
    .A2(_04913_),
    .ZN(_05871_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12571_ (.I0(_05869_),
    .I1(\mod.u_cpu.rf_ram.memory[15][0] ),
    .S(_05871_),
    .Z(_05872_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12572_ (.I(_05872_),
    .Z(_01003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12573_ (.I(_05709_),
    .Z(_05873_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12574_ (.I(_05873_),
    .Z(_05874_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12575_ (.I0(_05874_),
    .I1(\mod.u_cpu.rf_ram.memory[15][1] ),
    .S(_05871_),
    .Z(_05875_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12576_ (.I(_05875_),
    .Z(_01004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12577_ (.A1(_05428_),
    .A2(_05374_),
    .ZN(_05876_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12578_ (.I0(_05869_),
    .I1(\mod.u_cpu.rf_ram.memory[158][0] ),
    .S(_05876_),
    .Z(_05877_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12579_ (.I(_05877_),
    .Z(_01005_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12580_ (.I0(_05874_),
    .I1(\mod.u_cpu.rf_ram.memory[158][1] ),
    .S(_05876_),
    .Z(_05878_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12581_ (.I(_05878_),
    .Z(_01006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12582_ (.A1(_05515_),
    .A2(_05374_),
    .ZN(_05879_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12583_ (.I0(_05869_),
    .I1(\mod.u_cpu.rf_ram.memory[157][0] ),
    .S(_05879_),
    .Z(_05880_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12584_ (.I(_05880_),
    .Z(_01007_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12585_ (.I0(_05874_),
    .I1(\mod.u_cpu.rf_ram.memory[157][1] ),
    .S(_05879_),
    .Z(_05881_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12586_ (.I(_05881_),
    .Z(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12587_ (.I(_05373_),
    .Z(_05882_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12588_ (.A1(_05443_),
    .A2(_05882_),
    .ZN(_05883_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12589_ (.I0(_05869_),
    .I1(\mod.u_cpu.rf_ram.memory[156][0] ),
    .S(_05883_),
    .Z(_05884_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12590_ (.I(_05884_),
    .Z(_01009_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12591_ (.I0(_05874_),
    .I1(\mod.u_cpu.rf_ram.memory[156][1] ),
    .S(_05883_),
    .Z(_05885_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12592_ (.I(_05885_),
    .Z(_01010_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12593_ (.I(_05694_),
    .Z(_05886_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12594_ (.I(_05886_),
    .Z(_05887_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12595_ (.I(_03789_),
    .Z(_05888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12596_ (.A1(_05888_),
    .A2(_05882_),
    .ZN(_05889_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12597_ (.I0(_05887_),
    .I1(\mod.u_cpu.rf_ram.memory[155][0] ),
    .S(_05889_),
    .Z(_05890_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12598_ (.I(_05890_),
    .Z(_01011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12599_ (.I(_05873_),
    .Z(_05891_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12600_ (.I0(_05891_),
    .I1(\mod.u_cpu.rf_ram.memory[155][1] ),
    .S(_05889_),
    .Z(_05892_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12601_ (.I(_05892_),
    .Z(_01012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12602_ (.A1(_03796_),
    .A2(_05882_),
    .ZN(_05893_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12603_ (.I0(_05887_),
    .I1(\mod.u_cpu.rf_ram.memory[154][0] ),
    .S(_05893_),
    .Z(_05894_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12604_ (.I(_05894_),
    .Z(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12605_ (.I0(_05891_),
    .I1(\mod.u_cpu.rf_ram.memory[154][1] ),
    .S(_05893_),
    .Z(_05895_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12606_ (.I(_05895_),
    .Z(_01014_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12607_ (.I(_04024_),
    .Z(_05896_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12608_ (.A1(_05896_),
    .A2(_05882_),
    .ZN(_05897_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12609_ (.I0(_05887_),
    .I1(\mod.u_cpu.rf_ram.memory[153][0] ),
    .S(_05897_),
    .Z(_05898_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12610_ (.I(_05898_),
    .Z(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12611_ (.I0(_05891_),
    .I1(\mod.u_cpu.rf_ram.memory[153][1] ),
    .S(_05897_),
    .Z(_05899_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12612_ (.I(_05899_),
    .Z(_01016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12613_ (.I(_05373_),
    .Z(_05900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12614_ (.A1(_05283_),
    .A2(_05900_),
    .ZN(_05901_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12615_ (.I0(_05887_),
    .I1(\mod.u_cpu.rf_ram.memory[152][0] ),
    .S(_05901_),
    .Z(_05902_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12616_ (.I(_05902_),
    .Z(_01017_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12617_ (.I0(_05891_),
    .I1(\mod.u_cpu.rf_ram.memory[152][1] ),
    .S(_05901_),
    .Z(_05903_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12618_ (.I(_05903_),
    .Z(_01018_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12619_ (.I(_05886_),
    .Z(_05904_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12620_ (.A1(_03879_),
    .A2(_05900_),
    .ZN(_05905_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12621_ (.I0(_05904_),
    .I1(\mod.u_cpu.rf_ram.memory[151][0] ),
    .S(_05905_),
    .Z(_05906_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12622_ (.I(_05906_),
    .Z(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12623_ (.I(_05873_),
    .Z(_05907_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12624_ (.I0(_05907_),
    .I1(\mod.u_cpu.rf_ram.memory[151][1] ),
    .S(_05905_),
    .Z(_05908_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12625_ (.I(_05908_),
    .Z(_01020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12626_ (.A1(_05494_),
    .A2(_05900_),
    .ZN(_05909_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12627_ (.I0(_05904_),
    .I1(\mod.u_cpu.rf_ram.memory[150][0] ),
    .S(_05909_),
    .Z(_05910_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12628_ (.I(_05910_),
    .Z(_01021_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12629_ (.I0(_05907_),
    .I1(\mod.u_cpu.rf_ram.memory[150][1] ),
    .S(_05909_),
    .Z(_05911_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12630_ (.I(_05911_),
    .Z(_01022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12631_ (.A1(_05870_),
    .A2(_03886_),
    .ZN(_05912_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12632_ (.I0(_05904_),
    .I1(\mod.u_cpu.rf_ram.memory[14][0] ),
    .S(_05912_),
    .Z(_05913_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12633_ (.I(_05913_),
    .Z(_01023_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12634_ (.I0(_05907_),
    .I1(\mod.u_cpu.rf_ram.memory[14][1] ),
    .S(_05912_),
    .Z(_05914_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12635_ (.I(_05914_),
    .Z(_01024_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12636_ (.A1(_05535_),
    .A2(_05900_),
    .ZN(_05915_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12637_ (.I0(_05904_),
    .I1(\mod.u_cpu.rf_ram.memory[148][0] ),
    .S(_05915_),
    .Z(_05916_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12638_ (.I(_05916_),
    .Z(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12639_ (.I0(_05907_),
    .I1(\mod.u_cpu.rf_ram.memory[148][1] ),
    .S(_05915_),
    .Z(_05917_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12640_ (.I(_05917_),
    .Z(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12641_ (.I(_05886_),
    .Z(_05918_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12642_ (.I(_05372_),
    .Z(_05919_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12643_ (.I(_05919_),
    .Z(_05920_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12644_ (.A1(_05732_),
    .A2(_05920_),
    .ZN(_05921_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12645_ (.I0(_05918_),
    .I1(\mod.u_cpu.rf_ram.memory[147][0] ),
    .S(_05921_),
    .Z(_05922_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12646_ (.I(_05922_),
    .Z(_01027_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12647_ (.I(_05873_),
    .Z(_05923_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12648_ (.I0(_05923_),
    .I1(\mod.u_cpu.rf_ram.memory[147][1] ),
    .S(_05921_),
    .Z(_05924_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12649_ (.I(_05924_),
    .Z(_01028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12650_ (.A1(_05293_),
    .A2(_05920_),
    .ZN(_05925_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12651_ (.I0(_05918_),
    .I1(\mod.u_cpu.rf_ram.memory[146][0] ),
    .S(_05925_),
    .Z(_05926_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12652_ (.I(_05926_),
    .Z(_01029_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12653_ (.I0(_05923_),
    .I1(\mod.u_cpu.rf_ram.memory[146][1] ),
    .S(_05925_),
    .Z(_05927_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12654_ (.I(_05927_),
    .Z(_01030_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12655_ (.A1(_05742_),
    .A2(_05920_),
    .ZN(_05928_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12656_ (.I0(_05918_),
    .I1(\mod.u_cpu.rf_ram.memory[145][0] ),
    .S(_05928_),
    .Z(_05929_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12657_ (.I(_05929_),
    .Z(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12658_ (.I0(_05923_),
    .I1(\mod.u_cpu.rf_ram.memory[145][1] ),
    .S(_05928_),
    .Z(_05930_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12659_ (.I(_05930_),
    .Z(_01032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12660_ (.A1(_05300_),
    .A2(_05920_),
    .ZN(_05931_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12661_ (.I0(_05918_),
    .I1(\mod.u_cpu.rf_ram.memory[144][0] ),
    .S(_05931_),
    .Z(_05932_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12662_ (.I(_05932_),
    .Z(_01033_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12663_ (.I0(_05923_),
    .I1(\mod.u_cpu.rf_ram.memory[144][1] ),
    .S(_05931_),
    .Z(_05933_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12664_ (.I(_05933_),
    .Z(_01034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12665_ (.I(_05886_),
    .Z(_05934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12666_ (.A1(_05896_),
    .A2(_05721_),
    .ZN(_05935_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12667_ (.I0(_05934_),
    .I1(\mod.u_cpu.rf_ram.memory[121][0] ),
    .S(_05935_),
    .Z(_05936_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12668_ (.I(_05936_),
    .Z(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12669_ (.I(_05709_),
    .Z(_05937_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12670_ (.I(_05937_),
    .Z(_05938_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12671_ (.I0(_05938_),
    .I1(\mod.u_cpu.rf_ram.memory[121][1] ),
    .S(_05935_),
    .Z(_05939_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12672_ (.I(_05939_),
    .Z(_01036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12673_ (.I(_05919_),
    .Z(_05940_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12674_ (.A1(_04913_),
    .A2(_05940_),
    .ZN(_05941_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12675_ (.I0(_05934_),
    .I1(\mod.u_cpu.rf_ram.memory[143][0] ),
    .S(_05941_),
    .Z(_05942_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12676_ (.I(_05942_),
    .Z(_01037_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12677_ (.I0(_05938_),
    .I1(\mod.u_cpu.rf_ram.memory[143][1] ),
    .S(_05941_),
    .Z(_05943_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12678_ (.I(_05943_),
    .Z(_01038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12679_ (.A1(_05312_),
    .A2(_05940_),
    .ZN(_05944_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12680_ (.I0(_05934_),
    .I1(\mod.u_cpu.rf_ram.memory[142][0] ),
    .S(_05944_),
    .Z(_05945_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12681_ (.I(_05945_),
    .Z(_01039_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12682_ (.I0(_05938_),
    .I1(\mod.u_cpu.rf_ram.memory[142][1] ),
    .S(_05944_),
    .Z(_05946_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12683_ (.I(_05946_),
    .Z(_01040_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12684_ (.A1(_03895_),
    .A2(_05589_),
    .ZN(_05947_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12685_ (.I(_03944_),
    .Z(_05948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12686_ (.A1(_05948_),
    .A2(_05947_),
    .ZN(_05949_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12687_ (.A1(_02370_),
    .A2(_05947_),
    .B(_05949_),
    .ZN(_01041_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12688_ (.I(_03734_),
    .Z(_05950_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12689_ (.I0(\mod.u_cpu.rf_ram.memory[77][1] ),
    .I1(_05950_),
    .S(_05947_),
    .Z(_05951_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12690_ (.I(_05951_),
    .Z(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _12691_ (.A1(_03723_),
    .A2(_05319_),
    .ZN(_05952_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12692_ (.A1(_04643_),
    .A2(_05952_),
    .ZN(_05953_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12693_ (.I0(\mod.u_cpu.rf_ram.memory[141][0] ),
    .I1(_05622_),
    .S(_05953_),
    .Z(_05954_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12694_ (.I(_05954_),
    .Z(_01043_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12695_ (.I0(\mod.u_cpu.rf_ram.memory[141][1] ),
    .I1(_05950_),
    .S(_05953_),
    .Z(_05955_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12696_ (.I(_05955_),
    .Z(_01044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12697_ (.A1(_03904_),
    .A2(_05940_),
    .ZN(_05956_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12698_ (.I0(_05934_),
    .I1(\mod.u_cpu.rf_ram.memory[140][0] ),
    .S(_05956_),
    .Z(_05957_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12699_ (.I(_05957_),
    .Z(_01045_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12700_ (.I0(_05938_),
    .I1(\mod.u_cpu.rf_ram.memory[140][1] ),
    .S(_05956_),
    .Z(_05958_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12701_ (.I(_05958_),
    .Z(_01046_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12702_ (.A1(_03728_),
    .A2(_04643_),
    .ZN(_05959_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12703_ (.I0(\mod.u_cpu.rf_ram.memory[13][0] ),
    .I1(_05622_),
    .S(_05959_),
    .Z(_05960_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12704_ (.I(_05960_),
    .Z(_01047_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12705_ (.I0(\mod.u_cpu.rf_ram.memory[13][1] ),
    .I1(_05950_),
    .S(_05959_),
    .Z(_05961_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12706_ (.I(_05961_),
    .Z(_01048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12707_ (.I(_05694_),
    .Z(_05962_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12708_ (.I(_05962_),
    .Z(_05963_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12709_ (.A1(_05870_),
    .A2(_04668_),
    .ZN(_05964_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12710_ (.I0(_05963_),
    .I1(\mod.u_cpu.rf_ram.memory[7][0] ),
    .S(_05964_),
    .Z(_05965_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12711_ (.I(_05965_),
    .Z(_01049_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12712_ (.I(_05937_),
    .Z(_05966_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12713_ (.I0(_05966_),
    .I1(\mod.u_cpu.rf_ram.memory[7][1] ),
    .S(_05964_),
    .Z(_05967_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12714_ (.I(_05967_),
    .Z(_01050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12715_ (.A1(_03918_),
    .A2(_05940_),
    .ZN(_05968_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12716_ (.I0(_05963_),
    .I1(\mod.u_cpu.rf_ram.memory[138][0] ),
    .S(_05968_),
    .Z(_05969_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12717_ (.I(_05969_),
    .Z(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12718_ (.I0(_05966_),
    .I1(\mod.u_cpu.rf_ram.memory[138][1] ),
    .S(_05968_),
    .Z(_05970_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12719_ (.I(_05970_),
    .Z(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12720_ (.I(_03698_),
    .Z(_05971_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12721_ (.A1(_05588_),
    .A2(_05952_),
    .ZN(_05972_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12722_ (.I0(\mod.u_cpu.rf_ram.memory[137][0] ),
    .I1(_05971_),
    .S(_05972_),
    .Z(_05973_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12723_ (.I(_05973_),
    .Z(_01053_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12724_ (.I0(\mod.u_cpu.rf_ram.memory[137][1] ),
    .I1(_05950_),
    .S(_05972_),
    .Z(_05974_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12725_ (.I(_05974_),
    .Z(_01054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12726_ (.A1(_03885_),
    .A2(_05576_),
    .ZN(_05975_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12727_ (.I0(_05963_),
    .I1(\mod.u_cpu.rf_ram.memory[78][0] ),
    .S(_05975_),
    .Z(_05976_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12728_ (.I(_05976_),
    .Z(_01055_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12729_ (.I0(_05966_),
    .I1(\mod.u_cpu.rf_ram.memory[78][1] ),
    .S(_05975_),
    .Z(_05977_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12730_ (.I(_05977_),
    .Z(_01056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12731_ (.I(_05919_),
    .Z(_05978_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12732_ (.A1(_03932_),
    .A2(_05978_),
    .ZN(_05979_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12733_ (.I0(_05963_),
    .I1(\mod.u_cpu.rf_ram.memory[136][0] ),
    .S(_05979_),
    .Z(_05980_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12734_ (.I(_05980_),
    .Z(_01057_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12735_ (.I0(_05966_),
    .I1(\mod.u_cpu.rf_ram.memory[136][1] ),
    .S(_05979_),
    .Z(_05981_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12736_ (.I(_05981_),
    .Z(_01058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12737_ (.A1(_03865_),
    .A2(_05552_),
    .ZN(_05982_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12738_ (.A1(_05843_),
    .A2(_05982_),
    .ZN(_05983_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12739_ (.A1(_02215_),
    .A2(_05982_),
    .B(_05983_),
    .ZN(_01059_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12740_ (.I(_05937_),
    .Z(_05984_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12741_ (.I0(_05984_),
    .I1(\mod.u_cpu.rf_ram.memory[209][1] ),
    .S(_05982_),
    .Z(_05985_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12742_ (.I(_05985_),
    .Z(_01060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12743_ (.A1(_03790_),
    .A2(_05552_),
    .ZN(_05986_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12744_ (.A1(_05843_),
    .A2(_05986_),
    .ZN(_05987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12745_ (.A1(_02199_),
    .A2(_05986_),
    .B(_05987_),
    .ZN(_01061_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12746_ (.I0(_05984_),
    .I1(\mod.u_cpu.rf_ram.memory[219][1] ),
    .S(_05986_),
    .Z(_05988_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12747_ (.I(_05988_),
    .Z(_01062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12748_ (.A1(_05395_),
    .A2(_05422_),
    .ZN(_05989_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12749_ (.A1(_05843_),
    .A2(_05989_),
    .ZN(_05990_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12750_ (.A1(_02162_),
    .A2(_05989_),
    .B(_05990_),
    .ZN(_01063_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12751_ (.I0(_05984_),
    .I1(\mod.u_cpu.rf_ram.memory[199][1] ),
    .S(_05989_),
    .Z(_05991_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12752_ (.I(_05991_),
    .Z(_01064_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12753_ (.I(_05962_),
    .Z(_05992_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12754_ (.A1(_03872_),
    .A2(_05576_),
    .ZN(_05993_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12755_ (.I0(_05992_),
    .I1(\mod.u_cpu.rf_ram.memory[80][0] ),
    .S(_05993_),
    .Z(_05994_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12756_ (.I(_05994_),
    .Z(_01065_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12757_ (.I0(_05984_),
    .I1(\mod.u_cpu.rf_ram.memory[80][1] ),
    .S(_05993_),
    .Z(_05995_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12758_ (.I(_05995_),
    .Z(_01066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12759_ (.A1(_04668_),
    .A2(_05978_),
    .ZN(_05996_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12760_ (.I0(_05992_),
    .I1(\mod.u_cpu.rf_ram.memory[135][0] ),
    .S(_05996_),
    .Z(_05997_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12761_ (.I(_05997_),
    .Z(_01067_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12762_ (.I(_05937_),
    .Z(_05998_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12763_ (.I0(_05998_),
    .I1(\mod.u_cpu.rf_ram.memory[135][1] ),
    .S(_05996_),
    .Z(_05999_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12764_ (.I(_05999_),
    .Z(_01068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12765_ (.A1(_03950_),
    .A2(_05978_),
    .ZN(_06000_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12766_ (.I0(_05992_),
    .I1(\mod.u_cpu.rf_ram.memory[134][0] ),
    .S(_06000_),
    .Z(_06001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12767_ (.I(_06001_),
    .Z(_01069_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12768_ (.I0(_05998_),
    .I1(\mod.u_cpu.rf_ram.memory[134][1] ),
    .S(_06000_),
    .Z(_06002_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12769_ (.I(_06002_),
    .Z(_01070_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12770_ (.A1(_04955_),
    .A2(_05952_),
    .ZN(_06003_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12771_ (.I0(\mod.u_cpu.rf_ram.memory[133][0] ),
    .I1(_05971_),
    .S(_06003_),
    .Z(_06004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12772_ (.I(_06004_),
    .Z(_01071_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12773_ (.I(_03734_),
    .Z(_06005_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12774_ (.I0(\mod.u_cpu.rf_ram.memory[133][1] ),
    .I1(_06005_),
    .S(_06003_),
    .Z(_06006_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12775_ (.I(_06006_),
    .Z(_01072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12776_ (.A1(_03960_),
    .A2(_05978_),
    .ZN(_06007_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12777_ (.I0(_05992_),
    .I1(\mod.u_cpu.rf_ram.memory[132][0] ),
    .S(_06007_),
    .Z(_06008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12778_ (.I(_06008_),
    .Z(_01073_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12779_ (.I0(_05998_),
    .I1(\mod.u_cpu.rf_ram.memory[132][1] ),
    .S(_06007_),
    .Z(_06009_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12780_ (.I(_06009_),
    .Z(_01074_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12781_ (.I(_05962_),
    .Z(_06010_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12782_ (.I(_05919_),
    .Z(_06011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12783_ (.A1(_05649_),
    .A2(_06011_),
    .ZN(_06012_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12784_ (.I0(_06010_),
    .I1(\mod.u_cpu.rf_ram.memory[131][0] ),
    .S(_06012_),
    .Z(_06013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12785_ (.I(_06013_),
    .Z(_01075_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12786_ (.I0(_05998_),
    .I1(\mod.u_cpu.rf_ram.memory[131][1] ),
    .S(_06012_),
    .Z(_06014_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12787_ (.I(_06014_),
    .Z(_01076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12788_ (.A1(_03974_),
    .A2(_06011_),
    .ZN(_06015_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12789_ (.I0(_06010_),
    .I1(\mod.u_cpu.rf_ram.memory[130][0] ),
    .S(_06015_),
    .Z(_06016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12790_ (.I(_06016_),
    .Z(_01077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12791_ (.I(_05105_),
    .Z(_06017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12792_ (.I(_06017_),
    .Z(_06018_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12793_ (.I(_06018_),
    .Z(_06019_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12794_ (.I0(_06019_),
    .I1(\mod.u_cpu.rf_ram.memory[130][1] ),
    .S(_06015_),
    .Z(_06020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12795_ (.I(_06020_),
    .Z(_01078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12796_ (.A1(_05870_),
    .A2(_03905_),
    .ZN(_06021_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12797_ (.I0(_06010_),
    .I1(\mod.u_cpu.rf_ram.memory[12][0] ),
    .S(_06021_),
    .Z(_06022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12798_ (.I(_06022_),
    .Z(_01079_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12799_ (.I0(_06019_),
    .I1(\mod.u_cpu.rf_ram.memory[12][1] ),
    .S(_06021_),
    .Z(_06023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12800_ (.I(_06023_),
    .Z(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12801_ (.A1(_03985_),
    .A2(_06011_),
    .ZN(_06024_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12802_ (.I0(_06010_),
    .I1(\mod.u_cpu.rf_ram.memory[128][0] ),
    .S(_06024_),
    .Z(_06025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12803_ (.I(_06025_),
    .Z(_01081_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12804_ (.I0(_06019_),
    .I1(\mod.u_cpu.rf_ram.memory[128][1] ),
    .S(_06024_),
    .Z(_06026_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12805_ (.I(_06026_),
    .Z(_01082_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12806_ (.A1(_05226_),
    .A2(_05320_),
    .ZN(_06027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12807_ (.A1(_05948_),
    .A2(_06027_),
    .ZN(_06028_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12808_ (.A1(_02234_),
    .A2(_06027_),
    .B(_06028_),
    .ZN(_01083_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12809_ (.I0(\mod.u_cpu.rf_ram.memory[229][1] ),
    .I1(_06005_),
    .S(_06027_),
    .Z(_06029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12810_ (.I(_06029_),
    .Z(_01084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12811_ (.I(_05630_),
    .Z(_06030_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12812_ (.A1(_04844_),
    .A2(_06030_),
    .ZN(_06031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12813_ (.I(_03774_),
    .Z(_06032_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12814_ (.A1(_06032_),
    .A2(_06031_),
    .ZN(_06033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12815_ (.A1(_02317_),
    .A2(_06031_),
    .B(_06033_),
    .ZN(_01085_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12816_ (.I0(_06019_),
    .I1(\mod.u_cpu.rf_ram.memory[127][1] ),
    .S(_06031_),
    .Z(_06034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12817_ (.I(_06034_),
    .Z(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12818_ (.I(_05962_),
    .Z(_06035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12819_ (.A1(_03751_),
    .A2(_05721_),
    .ZN(_06036_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12820_ (.I0(_06035_),
    .I1(\mod.u_cpu.rf_ram.memory[126][0] ),
    .S(_06036_),
    .Z(_06037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12821_ (.I(_06037_),
    .Z(_01087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12822_ (.I(_06018_),
    .Z(_06038_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12823_ (.I0(_06038_),
    .I1(\mod.u_cpu.rf_ram.memory[126][1] ),
    .S(_06036_),
    .Z(_06039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12824_ (.I(_06039_),
    .Z(_01088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12825_ (.A1(_03770_),
    .A2(_06030_),
    .ZN(_06040_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12826_ (.A1(_06032_),
    .A2(_06040_),
    .ZN(_06041_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12827_ (.A1(_02313_),
    .A2(_06040_),
    .B(_06041_),
    .ZN(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12828_ (.I0(_06038_),
    .I1(\mod.u_cpu.rf_ram.memory[125][1] ),
    .S(_06040_),
    .Z(_06042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12829_ (.I(_06042_),
    .Z(_01090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12830_ (.A1(_03781_),
    .A2(_05721_),
    .ZN(_06043_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12831_ (.I0(_06035_),
    .I1(\mod.u_cpu.rf_ram.memory[124][0] ),
    .S(_06043_),
    .Z(_06044_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12832_ (.I(_06044_),
    .Z(_01091_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12833_ (.I0(_06038_),
    .I1(\mod.u_cpu.rf_ram.memory[124][1] ),
    .S(_06043_),
    .Z(_06045_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12834_ (.I(_06045_),
    .Z(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12835_ (.I(net5),
    .Z(_06046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12836_ (.I(_06046_),
    .Z(_06047_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12837_ (.A1(_06047_),
    .A2(_05788_),
    .ZN(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12838_ (.I(_05720_),
    .Z(_06048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12839_ (.A1(_05888_),
    .A2(_06048_),
    .ZN(_06049_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12840_ (.I0(_06035_),
    .I1(\mod.u_cpu.rf_ram.memory[123][0] ),
    .S(_06049_),
    .Z(_06050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12841_ (.I(_06050_),
    .Z(_01094_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12842_ (.I0(_06038_),
    .I1(\mod.u_cpu.rf_ram.memory[123][1] ),
    .S(_06049_),
    .Z(_06051_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12843_ (.I(_06051_),
    .Z(_01095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12844_ (.A1(_05788_),
    .A2(_05803_),
    .ZN(_06052_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12845_ (.A1(_01478_),
    .A2(_06052_),
    .ZN(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12846_ (.A1(_03743_),
    .A2(_06052_),
    .ZN(_01097_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12847_ (.A1(_02080_),
    .A2(_03742_),
    .Z(_06053_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12848_ (.A1(_06052_),
    .A2(_06053_),
    .ZN(_01098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12849_ (.A1(_02523_),
    .A2(_03742_),
    .ZN(_06054_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _12850_ (.A1(_02505_),
    .A2(_06054_),
    .Z(_06055_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12851_ (.A1(_06052_),
    .A2(_06055_),
    .ZN(_01099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12852_ (.I(_03398_),
    .Z(_06056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12853_ (.I(_06056_),
    .Z(_06057_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12854_ (.A1(_06057_),
    .A2(\mod.u_cpu.rf_ram_if.rreq_r ),
    .Z(_06058_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12855_ (.I(_06058_),
    .Z(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12856_ (.I(\mod.u_cpu.rf_ram.rdata[1] ),
    .ZN(_06059_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _12857_ (.A1(_01464_),
    .A2(\mod.u_cpu.rf_ram.regzero ),
    .A3(_06059_),
    .ZN(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12858_ (.I(\mod.u_cpu.rf_ram_if.rdata1 ),
    .ZN(_06060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12859_ (.A1(\mod.u_cpu.rf_ram_if.rtrig1 ),
    .A2(\mod.u_cpu.rf_ram.rdata[1] ),
    .ZN(_06061_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _12860_ (.A1(_06060_),
    .A2(\mod.u_cpu.rf_ram_if.rtrig1 ),
    .B1(_06061_),
    .B2(\mod.u_cpu.rf_ram.regzero ),
    .ZN(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12861_ (.I(_03338_),
    .Z(_06062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12862_ (.I(_06062_),
    .Z(_06063_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12863_ (.I(_05786_),
    .Z(_06064_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12864_ (.I(_06064_),
    .Z(_06065_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12865_ (.A1(_06063_),
    .A2(_06065_),
    .ZN(_06066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12866_ (.A1(\mod.u_cpu.cpu.state.ibus_cyc ),
    .A2(_06066_),
    .B(_06046_),
    .ZN(_06067_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12867_ (.A1(_03677_),
    .A2(_06066_),
    .B(_06067_),
    .ZN(_01103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12868_ (.A1(_05896_),
    .A2(_04687_),
    .ZN(_06068_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12869_ (.I0(_06035_),
    .I1(\mod.u_cpu.rf_ram.memory[409][0] ),
    .S(_06068_),
    .Z(_06069_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12870_ (.I(_06069_),
    .Z(_01104_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12871_ (.I(_06018_),
    .Z(_06070_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12872_ (.I0(_06070_),
    .I1(\mod.u_cpu.rf_ram.memory[409][1] ),
    .S(_06068_),
    .Z(_06071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12873_ (.I(_06071_),
    .Z(_01105_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12874_ (.I(_03923_),
    .Z(_06072_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12875_ (.I(_06072_),
    .Z(_06073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12876_ (.A1(_05494_),
    .A2(_05263_),
    .ZN(_06074_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12877_ (.I0(_06073_),
    .I1(\mod.u_cpu.rf_ram.memory[246][0] ),
    .S(_06074_),
    .Z(_06075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12878_ (.I(_06075_),
    .Z(_01106_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12879_ (.I0(_06070_),
    .I1(\mod.u_cpu.rf_ram.memory[246][1] ),
    .S(_06074_),
    .Z(_06076_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12880_ (.I(_06076_),
    .Z(_01107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12881_ (.A1(_03968_),
    .A2(_06048_),
    .ZN(_06077_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12882_ (.I0(_06073_),
    .I1(\mod.u_cpu.rf_ram.memory[99][0] ),
    .S(_06077_),
    .Z(_06078_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12883_ (.I(_06078_),
    .Z(_01108_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12884_ (.I0(_06070_),
    .I1(\mod.u_cpu.rf_ram.memory[99][1] ),
    .S(_06077_),
    .Z(_06079_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12885_ (.I(_06079_),
    .Z(_01109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12886_ (.I(_05396_),
    .Z(_06080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12887_ (.A1(_05896_),
    .A2(_06080_),
    .ZN(_06081_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12888_ (.I0(_06073_),
    .I1(\mod.u_cpu.rf_ram.memory[89][0] ),
    .S(_06081_),
    .Z(_06082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12889_ (.I(_06082_),
    .Z(_01110_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12890_ (.I0(_06070_),
    .I1(\mod.u_cpu.rf_ram.memory[89][1] ),
    .S(_06081_),
    .Z(_06083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12891_ (.I(_06083_),
    .Z(_01111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12892_ (.A1(_03974_),
    .A2(_06048_),
    .ZN(_06084_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12893_ (.I0(_06073_),
    .I1(\mod.u_cpu.rf_ram.memory[98][0] ),
    .S(_06084_),
    .Z(_06085_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12894_ (.I(_06085_),
    .Z(_01112_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12895_ (.I(_06018_),
    .Z(_06086_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12896_ (.I0(_06086_),
    .I1(\mod.u_cpu.rf_ram.memory[98][1] ),
    .S(_06084_),
    .Z(_06087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12897_ (.I(_06087_),
    .Z(_01113_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12898_ (.I(_06072_),
    .Z(_06088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12899_ (.A1(_03985_),
    .A2(_06048_),
    .ZN(_06089_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12900_ (.I0(_06088_),
    .I1(\mod.u_cpu.rf_ram.memory[96][0] ),
    .S(_06089_),
    .Z(_06090_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12901_ (.I(_06090_),
    .Z(_01114_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12902_ (.I0(_06086_),
    .I1(\mod.u_cpu.rf_ram.memory[96][1] ),
    .S(_06089_),
    .Z(_06091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12903_ (.I(_06091_),
    .Z(_01115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12904_ (.I(_05720_),
    .Z(_06092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12905_ (.A1(_05657_),
    .A2(_06092_),
    .ZN(_06093_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12906_ (.I0(_06088_),
    .I1(\mod.u_cpu.rf_ram.memory[97][0] ),
    .S(_06093_),
    .Z(_06094_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12907_ (.I(_06094_),
    .Z(_01116_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12908_ (.I0(_06086_),
    .I1(\mod.u_cpu.rf_ram.memory[97][1] ),
    .S(_06093_),
    .Z(_06095_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12909_ (.I(_06095_),
    .Z(_01117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12910_ (.A1(_04913_),
    .A2(_04570_),
    .ZN(_06096_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12911_ (.I0(_06088_),
    .I1(\mod.u_cpu.rf_ram.memory[399][0] ),
    .S(_06096_),
    .Z(_06097_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12912_ (.I(_06097_),
    .Z(_01118_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12913_ (.I0(_06086_),
    .I1(\mod.u_cpu.rf_ram.memory[399][1] ),
    .S(_06096_),
    .Z(_06098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12914_ (.I(_06098_),
    .Z(_01119_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _12915_ (.A1(_04955_),
    .A2(_04644_),
    .ZN(_06099_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12916_ (.I0(\mod.u_cpu.rf_ram.memory[389][0] ),
    .I1(_05971_),
    .S(_06099_),
    .Z(_06100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12917_ (.I(_06100_),
    .Z(_01120_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12918_ (.I0(\mod.u_cpu.rf_ram.memory[389][1] ),
    .I1(_06005_),
    .S(_06099_),
    .Z(_06101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12919_ (.I(_06101_),
    .Z(_01121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12920_ (.A1(_05888_),
    .A2(_04704_),
    .ZN(_06102_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12921_ (.I0(_06088_),
    .I1(\mod.u_cpu.rf_ram.memory[379][0] ),
    .S(_06102_),
    .Z(_06103_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12922_ (.I(_06103_),
    .Z(_01122_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12923_ (.I(_06017_),
    .Z(_06104_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12924_ (.I(_06104_),
    .Z(_06105_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12925_ (.I0(_06105_),
    .I1(\mod.u_cpu.rf_ram.memory[379][1] ),
    .S(_06102_),
    .Z(_06106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12926_ (.I(_06106_),
    .Z(_01123_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12927_ (.I(_06072_),
    .Z(_06107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12928_ (.A1(_05742_),
    .A2(_04704_),
    .ZN(_06108_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12929_ (.I0(_06107_),
    .I1(\mod.u_cpu.rf_ram.memory[369][0] ),
    .S(_06108_),
    .Z(_06109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12930_ (.I(_06109_),
    .Z(_01124_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12931_ (.I0(_06105_),
    .I1(\mod.u_cpu.rf_ram.memory[369][1] ),
    .S(_06108_),
    .Z(_06110_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12932_ (.I(_06110_),
    .Z(_01125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12933_ (.A1(_06062_),
    .A2(_03669_),
    .ZN(_06111_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12934_ (.A1(\mod.u_cpu.cpu.genblk3.csr.mie_mtie ),
    .A2(\mod.u_cpu.cpu.genblk3.csr.mstatus_mie ),
    .A3(\mod.timer_irq ),
    .ZN(_06112_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12935_ (.I(_01434_),
    .ZN(_06113_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _12936_ (.A1(\mod.u_cpu.cpu.genblk3.csr.timer_irq_r ),
    .A2(_06111_),
    .A3(_06112_),
    .B1(_06113_),
    .B2(_06063_),
    .ZN(_06114_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12937_ (.A1(_06057_),
    .A2(_06114_),
    .Z(_06115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12938_ (.I(_06115_),
    .Z(_01126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12939_ (.I(_05781_),
    .Z(_06116_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12940_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[14] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ),
    .S(_06116_),
    .Z(_06117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12941_ (.I(_06117_),
    .Z(_06118_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12942_ (.A1(_03500_),
    .A2(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ),
    .Z(_06119_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12943_ (.A1(_05784_),
    .A2(_03458_),
    .B(_06119_),
    .ZN(_06120_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12944_ (.A1(_06118_),
    .A2(_06120_),
    .ZN(_06121_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12945_ (.I(_03498_),
    .Z(_06122_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _12946_ (.I(\mod.u_arbiter.i_wb_cpu_rdt[0] ),
    .ZN(_06123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12947_ (.A1(_03500_),
    .A2(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ),
    .ZN(_06124_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12948_ (.A1(_06122_),
    .A2(_06123_),
    .B(_06124_),
    .ZN(_06125_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12949_ (.I(\mod.u_cpu.cpu.genblk1.align.ctrl_misal ),
    .Z(_06126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12950_ (.A1(_06116_),
    .A2(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ),
    .ZN(_06127_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12951_ (.A1(_06126_),
    .A2(_03424_),
    .B(_06127_),
    .ZN(_06128_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12952_ (.I(_06128_),
    .Z(_06129_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12953_ (.A1(_06125_),
    .A2(_06129_),
    .ZN(_06130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12954_ (.A1(_06125_),
    .A2(_06128_),
    .ZN(_06131_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12955_ (.I(_06131_),
    .ZN(_06132_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12956_ (.A1(_06121_),
    .A2(_06130_),
    .B(_06132_),
    .ZN(_06133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12957_ (.A1(_06064_),
    .A2(_06133_),
    .ZN(_06134_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12958_ (.I(_06134_),
    .Z(_06135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12959_ (.A1(\mod.u_arbiter.i_wb_cpu_ibus_adr[1] ),
    .A2(_05783_),
    .ZN(_06136_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _12960_ (.A1(\mod.u_arbiter.i_wb_cpu_ack ),
    .A2(_03399_),
    .A3(_06136_),
    .ZN(_06137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12961_ (.I(_06137_),
    .Z(_06138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12962_ (.I(_06138_),
    .Z(_06139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12963_ (.I(_06139_),
    .Z(_06140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12964_ (.A1(\mod.u_cpu.cpu.ctrl.i_iscomp ),
    .A2(_06140_),
    .ZN(_06141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12965_ (.A1(_06135_),
    .A2(_06141_),
    .ZN(_01127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12966_ (.I(_01425_),
    .Z(_06142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12967_ (.A1(_03338_),
    .A2(_03375_),
    .ZN(_06143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12968_ (.A1(_06142_),
    .A2(_06143_),
    .ZN(_06144_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12969_ (.A1(_03344_),
    .A2(_06144_),
    .ZN(_06145_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12970_ (.I(_03369_),
    .ZN(_06146_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12971_ (.A1(\mod.u_cpu.cpu.genblk3.csr.mstatus_mpie ),
    .A2(_06142_),
    .ZN(_06147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _12972_ (.A1(_06142_),
    .A2(_06146_),
    .B(_06147_),
    .C(_06145_),
    .ZN(_06148_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _12973_ (.A1(\mod.u_cpu.cpu.genblk3.csr.mstatus_mie ),
    .A2(_06145_),
    .B1(_06148_),
    .B2(_03353_),
    .ZN(_06149_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12974_ (.I(_06149_),
    .ZN(_01128_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _12975_ (.A1(_03389_),
    .A2(\mod.u_cpu.cpu.state.o_cnt[2] ),
    .Z(_06150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12976_ (.I(_06150_),
    .Z(_06151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12977_ (.I(_03269_),
    .Z(_06152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12978_ (.I(_03268_),
    .Z(_06153_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _12979_ (.A1(_01453_),
    .A2(_06152_),
    .A3(_06153_),
    .ZN(_06154_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _12980_ (.A1(\mod.u_cpu.cpu.decode.op22 ),
    .A2(_03343_),
    .A3(_06151_),
    .A4(_06154_),
    .Z(_06155_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12981_ (.A1(\mod.u_cpu.cpu.genblk3.csr.mie_mtie ),
    .A2(_06155_),
    .B(_06056_),
    .ZN(_06156_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12982_ (.A1(_06146_),
    .A2(_06155_),
    .B(_06156_),
    .ZN(_01129_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12983_ (.I0(\mod.u_cpu.cpu.genblk3.csr.mstatus_mie ),
    .I1(\mod.u_cpu.cpu.genblk3.csr.mstatus_mpie ),
    .S(_06143_),
    .Z(_06157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12984_ (.I(_06157_),
    .Z(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _12985_ (.A1(_06113_),
    .A2(_03370_),
    .ZN(_06158_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12986_ (.A1(_06063_),
    .A2(_03335_),
    .B(_03375_),
    .ZN(_06159_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12987_ (.I0(_06158_),
    .I1(\mod.u_cpu.cpu.genblk3.csr.mcause31 ),
    .S(_06159_),
    .Z(_06160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12988_ (.I(_06160_),
    .Z(_01131_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12989_ (.I(\mod.u_cpu.cpu.genblk3.csr.mcause3_0[1] ),
    .ZN(_06161_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _12990_ (.A1(_05780_),
    .A2(_06161_),
    .B(_03373_),
    .ZN(_06162_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _12991_ (.A1(_06062_),
    .A2(_03375_),
    .B1(_03337_),
    .B2(_03336_),
    .ZN(_06163_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _12992_ (.I(_06163_),
    .Z(_06164_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _12993_ (.I0(_06162_),
    .I1(\mod.u_cpu.cpu.genblk3.csr.mcause3_0[0] ),
    .S(_06164_),
    .Z(_06165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12994_ (.I(_06165_),
    .Z(_01132_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12995_ (.I(_03686_),
    .Z(_06166_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _12996_ (.I(\mod.u_cpu.cpu.genblk3.csr.mcause3_0[2] ),
    .ZN(_06167_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _12997_ (.A1(_06166_),
    .A2(_03404_),
    .B1(_06167_),
    .B2(_05780_),
    .C(_03373_),
    .ZN(_06168_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _12998_ (.A1(_06164_),
    .A2(_06168_),
    .ZN(_06169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _12999_ (.A1(_06161_),
    .A2(_06164_),
    .B(_06169_),
    .ZN(_01133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13000_ (.A1(_06113_),
    .A2(_06166_),
    .ZN(_06170_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _13001_ (.A1(\mod.u_cpu.cpu.genblk3.csr.mcause3_0[3] ),
    .A2(_03353_),
    .B(_06163_),
    .C(_06170_),
    .ZN(_06171_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13002_ (.A1(_06167_),
    .A2(_06164_),
    .B(_06171_),
    .ZN(_01134_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13003_ (.A1(_01435_),
    .A2(_01420_),
    .A3(_01424_),
    .ZN(_06172_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13004_ (.A1(_01453_),
    .A2(_06172_),
    .B(_03370_),
    .ZN(_06173_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13005_ (.I0(_06173_),
    .I1(\mod.u_cpu.cpu.genblk3.csr.mcause3_0[3] ),
    .S(_06163_),
    .Z(_06174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13006_ (.I(_06174_),
    .Z(_01135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13007_ (.A1(_03828_),
    .A2(_06080_),
    .ZN(_06175_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13008_ (.I0(_06107_),
    .I1(\mod.u_cpu.rf_ram.memory[86][0] ),
    .S(_06175_),
    .Z(_06176_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13009_ (.I(_06176_),
    .Z(_01136_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13010_ (.I0(_06105_),
    .I1(\mod.u_cpu.rf_ram.memory[86][1] ),
    .S(_06175_),
    .Z(_06177_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13011_ (.I(_06177_),
    .Z(_01137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13012_ (.A1(_03837_),
    .A2(_06080_),
    .ZN(_06178_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13013_ (.I0(_06107_),
    .I1(\mod.u_cpu.rf_ram.memory[85][0] ),
    .S(_06178_),
    .Z(_06179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13014_ (.I(_06179_),
    .Z(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13015_ (.I0(_06105_),
    .I1(\mod.u_cpu.rf_ram.memory[85][1] ),
    .S(_06178_),
    .Z(_06180_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13016_ (.I(_06180_),
    .Z(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13017_ (.I(_04982_),
    .Z(_06181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13018_ (.A1(_06181_),
    .A2(_03919_),
    .ZN(_06182_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13019_ (.I0(_06107_),
    .I1(\mod.u_cpu.rf_ram.memory[10][0] ),
    .S(_06182_),
    .Z(_06183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13020_ (.I(_06183_),
    .Z(_01140_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13021_ (.I(_06104_),
    .Z(_06184_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13022_ (.I0(_06184_),
    .I1(\mod.u_cpu.rf_ram.memory[10][1] ),
    .S(_06182_),
    .Z(_06185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13023_ (.I(_06185_),
    .Z(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13024_ (.I(_06072_),
    .Z(_06186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13025_ (.A1(_05535_),
    .A2(_06080_),
    .ZN(_06187_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13026_ (.I0(_06186_),
    .I1(\mod.u_cpu.rf_ram.memory[84][0] ),
    .S(_06187_),
    .Z(_06188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13027_ (.I(_06188_),
    .Z(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13028_ (.I0(_06184_),
    .I1(\mod.u_cpu.rf_ram.memory[84][1] ),
    .S(_06187_),
    .Z(_06189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13029_ (.I(_06189_),
    .Z(_01143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13030_ (.A1(_03904_),
    .A2(_06092_),
    .ZN(_06190_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13031_ (.I0(_06186_),
    .I1(\mod.u_cpu.rf_ram.memory[108][0] ),
    .S(_06190_),
    .Z(_06191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13032_ (.I(_06191_),
    .Z(_01144_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13033_ (.I0(_06184_),
    .I1(\mod.u_cpu.rf_ram.memory[108][1] ),
    .S(_06190_),
    .Z(_06192_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13034_ (.I(_06192_),
    .Z(_01145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13035_ (.I(_05396_),
    .Z(_06193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13036_ (.A1(_05732_),
    .A2(_06193_),
    .ZN(_06194_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13037_ (.I0(_06186_),
    .I1(\mod.u_cpu.rf_ram.memory[83][0] ),
    .S(_06194_),
    .Z(_06195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13038_ (.I(_06195_),
    .Z(_01146_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13039_ (.I0(_06184_),
    .I1(\mod.u_cpu.rf_ram.memory[83][1] ),
    .S(_06194_),
    .Z(_06196_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13040_ (.I(_06196_),
    .Z(_01147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13041_ (.A1(_05606_),
    .A2(_06092_),
    .ZN(_06197_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13042_ (.I0(_06186_),
    .I1(\mod.u_cpu.rf_ram.memory[107][0] ),
    .S(_06197_),
    .Z(_06198_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13043_ (.I(_06198_),
    .Z(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13044_ (.I(_06104_),
    .Z(_06199_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13045_ (.I0(_06199_),
    .I1(\mod.u_cpu.rf_ram.memory[107][1] ),
    .S(_06197_),
    .Z(_06200_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13046_ (.I(_06200_),
    .Z(_01149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13047_ (.A1(_04067_),
    .A2(_05387_),
    .ZN(_06201_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13048_ (.A1(_06032_),
    .A2(_06201_),
    .ZN(_06202_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13049_ (.A1(_02373_),
    .A2(_06201_),
    .B(_06202_),
    .ZN(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13050_ (.I0(_06199_),
    .I1(\mod.u_cpu.rf_ram.memory[79][1] ),
    .S(_06201_),
    .Z(_06203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13051_ (.I(_06203_),
    .Z(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13052_ (.I(_03923_),
    .Z(_06204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13053_ (.I(_06204_),
    .Z(_06205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13054_ (.A1(_03858_),
    .A2(_06193_),
    .ZN(_06206_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13055_ (.I0(_06205_),
    .I1(\mod.u_cpu.rf_ram.memory[82][0] ),
    .S(_06206_),
    .Z(_06207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13056_ (.I(_06207_),
    .Z(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13057_ (.I0(_06199_),
    .I1(\mod.u_cpu.rf_ram.memory[82][1] ),
    .S(_06206_),
    .Z(_06208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13058_ (.I(_06208_),
    .Z(_01153_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _13059_ (.A1(_04107_),
    .A2(_05589_),
    .ZN(_06209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13060_ (.A1(_05948_),
    .A2(_06209_),
    .ZN(_06210_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13061_ (.A1(_02353_),
    .A2(_06209_),
    .B(_06210_),
    .ZN(_01154_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13062_ (.I0(\mod.u_cpu.rf_ram.memory[69][1] ),
    .I1(_06005_),
    .S(_06209_),
    .Z(_06211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13063_ (.I(_06211_),
    .Z(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13064_ (.A1(_03918_),
    .A2(_06092_),
    .ZN(_06212_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13065_ (.I0(_06205_),
    .I1(\mod.u_cpu.rf_ram.memory[106][0] ),
    .S(_06212_),
    .Z(_06213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13066_ (.I(_06213_),
    .Z(_01156_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13067_ (.I0(_06199_),
    .I1(\mod.u_cpu.rf_ram.memory[106][1] ),
    .S(_06212_),
    .Z(_06214_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13068_ (.I(_06214_),
    .Z(_01157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13069_ (.A1(_05742_),
    .A2(_06193_),
    .ZN(_06215_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13070_ (.I0(_06205_),
    .I1(\mod.u_cpu.rf_ram.memory[81][0] ),
    .S(_06215_),
    .Z(_06216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13071_ (.I(_06216_),
    .Z(_01158_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13072_ (.I(_06104_),
    .Z(_06217_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13073_ (.I0(_06217_),
    .I1(\mod.u_cpu.rf_ram.memory[81][1] ),
    .S(_06215_),
    .Z(_06218_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13074_ (.I(_06218_),
    .Z(_01159_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _13075_ (.A1(_03713_),
    .A2(_05640_),
    .ZN(_06219_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13076_ (.I0(\mod.u_cpu.rf_ram.memory[105][0] ),
    .I1(_05971_),
    .S(_06219_),
    .Z(_06220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13077_ (.I(_06220_),
    .Z(_01160_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13078_ (.I(_03734_),
    .Z(_06221_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13079_ (.I0(\mod.u_cpu.rf_ram.memory[105][1] ),
    .I1(_06221_),
    .S(_06219_),
    .Z(_06222_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13080_ (.I(_06222_),
    .Z(_01161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13081_ (.I(_05630_),
    .Z(_06223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13082_ (.A1(_03932_),
    .A2(_06223_),
    .ZN(_06224_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13083_ (.I0(_06205_),
    .I1(\mod.u_cpu.rf_ram.memory[104][0] ),
    .S(_06224_),
    .Z(_06225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13084_ (.I(_06225_),
    .Z(_01162_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13085_ (.I0(_06217_),
    .I1(\mod.u_cpu.rf_ram.memory[104][1] ),
    .S(_06224_),
    .Z(_06226_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13086_ (.I(_06226_),
    .Z(_01163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13087_ (.A1(_03941_),
    .A2(_06030_),
    .ZN(_06227_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13088_ (.A1(_06032_),
    .A2(_06227_),
    .ZN(_06228_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13089_ (.A1(_02287_),
    .A2(_06227_),
    .B(_06228_),
    .ZN(_01164_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13090_ (.I0(_06217_),
    .I1(\mod.u_cpu.rf_ram.memory[103][1] ),
    .S(_06227_),
    .Z(_06229_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13091_ (.I(_06229_),
    .Z(_01165_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13092_ (.I(_06204_),
    .Z(_06230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13093_ (.A1(_05888_),
    .A2(_03878_),
    .ZN(_06231_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13094_ (.I0(_06230_),
    .I1(\mod.u_cpu.rf_ram.memory[59][0] ),
    .S(_06231_),
    .Z(_06232_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13095_ (.I(_06232_),
    .Z(_01166_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13096_ (.I0(_06217_),
    .I1(\mod.u_cpu.rf_ram.memory[59][1] ),
    .S(_06231_),
    .Z(_06233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13097_ (.I(_06233_),
    .Z(_01167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13098_ (.A1(_03950_),
    .A2(_06223_),
    .ZN(_06234_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13099_ (.I0(_06230_),
    .I1(\mod.u_cpu.rf_ram.memory[102][0] ),
    .S(_06234_),
    .Z(_06235_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13100_ (.I(_06235_),
    .Z(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13101_ (.I(_06017_),
    .Z(_06236_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13102_ (.I(_06236_),
    .Z(_06237_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13103_ (.I0(_06237_),
    .I1(\mod.u_cpu.rf_ram.memory[102][1] ),
    .S(_06234_),
    .Z(_06238_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13104_ (.I(_06238_),
    .Z(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _13105_ (.A1(_04107_),
    .A2(_05640_),
    .ZN(_06239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13106_ (.A1(_05948_),
    .A2(_06239_),
    .ZN(_06240_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13107_ (.A1(_02284_),
    .A2(_06239_),
    .B(_06240_),
    .ZN(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13108_ (.I0(\mod.u_cpu.rf_ram.memory[101][1] ),
    .I1(_06221_),
    .S(_06239_),
    .Z(_06241_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13109_ (.I(_06241_),
    .Z(_01171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13110_ (.A1(_03960_),
    .A2(_06223_),
    .ZN(_06242_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13111_ (.I0(_06230_),
    .I1(\mod.u_cpu.rf_ram.memory[100][0] ),
    .S(_06242_),
    .Z(_06243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13112_ (.I(_06243_),
    .Z(_01172_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13113_ (.I0(_06237_),
    .I1(\mod.u_cpu.rf_ram.memory[100][1] ),
    .S(_06242_),
    .Z(_06244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13114_ (.I(_06244_),
    .Z(_01173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13115_ (.A1(_06181_),
    .A2(_03986_),
    .ZN(_06245_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13116_ (.I0(_06230_),
    .I1(\mod.u_cpu.rf_ram.memory[0][0] ),
    .S(_06245_),
    .Z(_06246_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13117_ (.I(_06246_),
    .Z(_01174_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13118_ (.I0(_06237_),
    .I1(\mod.u_cpu.rf_ram.memory[0][1] ),
    .S(_06245_),
    .Z(_06247_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13119_ (.I(_06247_),
    .Z(_01175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13120_ (.A1(_03941_),
    .A2(_04708_),
    .ZN(_06248_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13121_ (.I(_03774_),
    .Z(_06249_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13122_ (.A1(_06249_),
    .A2(_06248_),
    .ZN(_06250_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13123_ (.A1(_01906_),
    .A2(_06248_),
    .B(_06250_),
    .ZN(_01176_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13124_ (.I0(_06237_),
    .I1(\mod.u_cpu.rf_ram.memory[359][1] ),
    .S(_06248_),
    .Z(_06251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13125_ (.I(_06251_),
    .Z(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13126_ (.I(_05785_),
    .Z(_06252_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13127_ (.I(_06252_),
    .Z(_06253_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13128_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[16] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ),
    .S(_06253_),
    .Z(_06254_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13129_ (.I(_06254_),
    .Z(_01178_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13130_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[17] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ),
    .S(_06253_),
    .Z(_06255_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13131_ (.I(_06255_),
    .Z(_01179_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13132_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[18] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[2] ),
    .S(_06253_),
    .Z(_06256_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13133_ (.I(_06256_),
    .Z(_01180_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13134_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[19] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[3] ),
    .S(_06253_),
    .Z(_06257_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13135_ (.I(_06257_),
    .Z(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13136_ (.I(_06252_),
    .Z(_06258_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13137_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[20] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ),
    .S(_06258_),
    .Z(_06259_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13138_ (.I(_06259_),
    .Z(_01182_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13139_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[21] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ),
    .S(_06258_),
    .Z(_06260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13140_ (.I(_06260_),
    .Z(_01183_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13141_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[22] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ),
    .S(_06258_),
    .Z(_06261_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13142_ (.I(_06261_),
    .Z(_01184_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13143_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[23] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ),
    .S(_06258_),
    .Z(_06262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13144_ (.I(_06262_),
    .Z(_01185_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13145_ (.I(_06252_),
    .Z(_06263_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13146_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[24] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ),
    .S(_06263_),
    .Z(_06264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13147_ (.I(_06264_),
    .Z(_01186_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13148_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[25] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ),
    .S(_06263_),
    .Z(_06265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13149_ (.I(_06265_),
    .Z(_01187_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13150_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[26] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[10] ),
    .S(_06263_),
    .Z(_06266_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13151_ (.I(_06266_),
    .Z(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13152_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[27] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[11] ),
    .S(_06263_),
    .Z(_06267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13153_ (.I(_06267_),
    .Z(_01189_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13154_ (.I(_06252_),
    .Z(_06268_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13155_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[28] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ),
    .S(_06268_),
    .Z(_06269_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13156_ (.I(_06269_),
    .Z(_01190_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13157_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[29] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ),
    .S(_06268_),
    .Z(_06270_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13158_ (.I(_06270_),
    .Z(_01191_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13159_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[30] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ),
    .S(_06268_),
    .Z(_06271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13160_ (.I(_06271_),
    .Z(_01192_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13161_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[31] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ),
    .S(_06268_),
    .Z(_06272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13162_ (.I(_06272_),
    .Z(_01193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13163_ (.I(_06204_),
    .Z(_06273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13164_ (.A1(_05515_),
    .A2(_04969_),
    .ZN(_06274_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13165_ (.I0(_06273_),
    .I1(\mod.u_cpu.rf_ram.memory[349][0] ),
    .S(_06274_),
    .Z(_06275_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13166_ (.I(_06275_),
    .Z(_01194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13167_ (.I(_06236_),
    .Z(_06276_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13168_ (.I0(_06276_),
    .I1(\mod.u_cpu.rf_ram.memory[349][1] ),
    .S(_06274_),
    .Z(_06277_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13169_ (.I(_06277_),
    .Z(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13170_ (.A1(_03492_),
    .A2(_03412_),
    .A3(_03400_),
    .ZN(_06278_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13171_ (.A1(_03510_),
    .A2(_06278_),
    .Z(_06279_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13172_ (.A1(_06047_),
    .A2(_06279_),
    .ZN(_01196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13173_ (.A1(\mod.u_cpu.cpu.bufreg.i_sh_signed ),
    .A2(_06140_),
    .ZN(_06280_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13174_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[10] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[10] ),
    .S(_05781_),
    .Z(_06281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13175_ (.I(_06281_),
    .Z(_06282_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13176_ (.I(_06282_),
    .Z(_06283_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13177_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[11] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[11] ),
    .S(_05781_),
    .Z(_06284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13178_ (.I(_06284_),
    .Z(_06285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13179_ (.A1(_06122_),
    .A2(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ),
    .ZN(_06286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13180_ (.A1(_05783_),
    .A2(\mod.u_arbiter.i_wb_cpu_rdt[12] ),
    .ZN(_06287_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13181_ (.A1(_06286_),
    .A2(_06287_),
    .Z(_06288_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13182_ (.I(_06288_),
    .Z(_06289_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13183_ (.A1(_03500_),
    .A2(\mod.u_arbiter.i_wb_cpu_rdt[5] ),
    .Z(_06290_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13184_ (.A1(_05783_),
    .A2(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ),
    .B(_06290_),
    .ZN(_06291_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13185_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[6] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ),
    .S(_06126_),
    .Z(_06292_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _13186_ (.I(_06292_),
    .ZN(_06293_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13187_ (.I(_06284_),
    .Z(_06294_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _13188_ (.A1(_06291_),
    .A2(_06293_),
    .A3(_06281_),
    .A4(_06294_),
    .ZN(_06295_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _13189_ (.A1(_06282_),
    .A2(_06289_),
    .B(_06295_),
    .C(_06285_),
    .ZN(_06296_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13190_ (.A1(_06116_),
    .A2(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ),
    .Z(_06297_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _13191_ (.A1(_05782_),
    .A2(_03456_),
    .B(_06297_),
    .ZN(_06298_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13192_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[15] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ),
    .S(_03499_),
    .Z(_06299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13193_ (.I(_06299_),
    .Z(_06300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13194_ (.A1(_06298_),
    .A2(_06300_),
    .ZN(_06301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13195_ (.A1(_06126_),
    .A2(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ),
    .ZN(_06302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13196_ (.A1(_05782_),
    .A2(\mod.u_arbiter.i_wb_cpu_rdt[13] ),
    .ZN(_06303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13197_ (.A1(_06302_),
    .A2(_06303_),
    .ZN(_06304_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _13198_ (.A1(_06301_),
    .A2(_06304_),
    .ZN(_06305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13199_ (.I(_06305_),
    .Z(_06306_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _13200_ (.A1(_06283_),
    .A2(_06285_),
    .B(_06296_),
    .C(_06306_),
    .ZN(_06307_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13201_ (.A1(_06302_),
    .A2(_06303_),
    .Z(_06308_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13202_ (.I(_06308_),
    .Z(_06309_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13203_ (.A1(_06118_),
    .A2(_06309_),
    .ZN(_06310_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13204_ (.I(_06310_),
    .Z(_06311_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13205_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[8] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ),
    .S(_03499_),
    .Z(_06312_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13206_ (.I(_06312_),
    .Z(_06313_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13207_ (.I(_06313_),
    .Z(_06314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13208_ (.A1(_06311_),
    .A2(_06314_),
    .ZN(_06315_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13209_ (.A1(_06117_),
    .A2(_06300_),
    .ZN(_06316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13210_ (.A1(_06309_),
    .A2(_06316_),
    .ZN(_06317_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13211_ (.I(_06317_),
    .Z(_06318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13212_ (.I(_06318_),
    .Z(_06319_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13213_ (.I(_06118_),
    .Z(_06320_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13214_ (.I(_06320_),
    .Z(_06321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13215_ (.A1(_06286_),
    .A2(_06287_),
    .ZN(_06322_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13216_ (.I(_06322_),
    .Z(_06323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13217_ (.A1(_06321_),
    .A2(_06323_),
    .ZN(_06324_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _13218_ (.A1(_06307_),
    .A2(_06315_),
    .A3(_06319_),
    .A4(_06324_),
    .ZN(_06325_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13219_ (.I(_06317_),
    .Z(_06326_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13220_ (.A1(_06122_),
    .A2(_06123_),
    .ZN(_06327_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13221_ (.A1(_03501_),
    .A2(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ),
    .B(_06327_),
    .ZN(_06328_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13222_ (.A1(_06328_),
    .A2(_06129_),
    .ZN(_06329_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13223_ (.I(_06329_),
    .Z(_06330_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13224_ (.A1(_06323_),
    .A2(_06326_),
    .B(_06330_),
    .ZN(_06331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13225_ (.I(_06331_),
    .Z(_06332_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13226_ (.A1(_06139_),
    .A2(_06332_),
    .ZN(_06333_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13227_ (.I(_03502_),
    .Z(_06334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13228_ (.I(_06334_),
    .Z(_06335_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13229_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[30] ),
    .I1(_03456_),
    .S(_06335_),
    .Z(_06336_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13230_ (.A1(_06137_),
    .A2(_06133_),
    .ZN(_06337_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13231_ (.I(_06337_),
    .Z(_06338_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13232_ (.I(_06338_),
    .Z(_06339_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13233_ (.A1(_06325_),
    .A2(_06333_),
    .B1(_06336_),
    .B2(_06339_),
    .ZN(_06340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13234_ (.A1(_06280_),
    .A2(_06340_),
    .ZN(_01197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13235_ (.A1(_03751_),
    .A2(_06193_),
    .ZN(_06341_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13236_ (.I0(_06273_),
    .I1(\mod.u_cpu.rf_ram.memory[94][0] ),
    .S(_06341_),
    .Z(_06342_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13237_ (.I(_06342_),
    .Z(_01198_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13238_ (.I0(_06276_),
    .I1(\mod.u_cpu.rf_ram.memory[94][1] ),
    .S(_06341_),
    .Z(_06343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13239_ (.I(_06343_),
    .Z(_01199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13240_ (.I(_05396_),
    .Z(_06344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13241_ (.A1(_03771_),
    .A2(_06344_),
    .ZN(_06345_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13242_ (.I0(_06273_),
    .I1(\mod.u_cpu.rf_ram.memory[93][0] ),
    .S(_06345_),
    .Z(_06346_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13243_ (.I(_06346_),
    .Z(_01200_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13244_ (.I0(_06276_),
    .I1(\mod.u_cpu.rf_ram.memory[93][1] ),
    .S(_06345_),
    .Z(_06347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13245_ (.I(_06347_),
    .Z(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13246_ (.A1(_03781_),
    .A2(_06344_),
    .ZN(_06348_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13247_ (.I0(_06273_),
    .I1(\mod.u_cpu.rf_ram.memory[92][0] ),
    .S(_06348_),
    .Z(_06349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13248_ (.I(_06349_),
    .Z(_01202_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13249_ (.I0(_06276_),
    .I1(\mod.u_cpu.rf_ram.memory[92][1] ),
    .S(_06348_),
    .Z(_06350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13250_ (.I(_06350_),
    .Z(_01203_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13251_ (.I(_06204_),
    .Z(_06351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13252_ (.A1(_04984_),
    .A2(_06344_),
    .ZN(_06352_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13253_ (.I0(_06351_),
    .I1(\mod.u_cpu.rf_ram.memory[95][0] ),
    .S(_06352_),
    .Z(_06353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13254_ (.I(_06353_),
    .Z(_01204_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13255_ (.I(_06236_),
    .Z(_06354_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13256_ (.I0(_06354_),
    .I1(\mod.u_cpu.rf_ram.memory[95][1] ),
    .S(_06352_),
    .Z(_06355_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13257_ (.I(_06355_),
    .Z(_01205_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13258_ (.A1(_03390_),
    .A2(_03672_),
    .ZN(_06356_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13259_ (.A1(_05787_),
    .A2(_06356_),
    .ZN(_06357_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13260_ (.I(_06357_),
    .Z(_06358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13261_ (.A1(_06126_),
    .A2(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ),
    .ZN(_06359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13262_ (.A1(_05782_),
    .A2(\mod.u_arbiter.i_wb_cpu_rdt[7] ),
    .ZN(_06360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13263_ (.A1(_06359_),
    .A2(_06360_),
    .ZN(_06361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13264_ (.I(_06361_),
    .Z(_06362_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13265_ (.I(_06362_),
    .Z(_06363_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13266_ (.I(_06361_),
    .Z(_06364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13267_ (.I(_06329_),
    .Z(_06365_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13268_ (.A1(_06318_),
    .A2(_06364_),
    .B(_06365_),
    .ZN(_06366_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13269_ (.I(_06298_),
    .Z(_06367_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13270_ (.I(_06120_),
    .Z(_06368_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13271_ (.A1(_06367_),
    .A2(_06368_),
    .ZN(_06369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13272_ (.I(_06369_),
    .Z(_06370_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13273_ (.I(_06322_),
    .Z(_06371_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13274_ (.I(_06371_),
    .Z(_06372_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13275_ (.A1(_06359_),
    .A2(_06360_),
    .Z(_06373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13276_ (.I(_06300_),
    .Z(_06374_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13277_ (.A1(_06321_),
    .A2(_06373_),
    .B(_06374_),
    .ZN(_06375_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _13278_ (.A1(_06306_),
    .A2(_06364_),
    .B1(_06370_),
    .B2(_06372_),
    .C(_06375_),
    .ZN(_06376_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13279_ (.I(_06116_),
    .Z(_06377_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13280_ (.A1(_06377_),
    .A2(_03424_),
    .ZN(_06378_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13281_ (.A1(_03501_),
    .A2(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ),
    .B(_06378_),
    .ZN(_06379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13282_ (.A1(_06328_),
    .A2(_06379_),
    .ZN(_06380_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13283_ (.I(_06380_),
    .Z(_06381_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13284_ (.I(_06368_),
    .Z(_06382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13285_ (.A1(_06367_),
    .A2(_06382_),
    .ZN(_06383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13286_ (.A1(_06291_),
    .A2(_06293_),
    .ZN(_06384_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13287_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[3] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[3] ),
    .S(_06377_),
    .Z(_06385_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13288_ (.A1(_06377_),
    .A2(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[2] ),
    .ZN(_06386_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13289_ (.A1(_03501_),
    .A2(_03428_),
    .B(_06386_),
    .ZN(_06387_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13290_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[4] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ),
    .S(_06122_),
    .Z(_06388_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _13291_ (.A1(_06384_),
    .A2(_06385_),
    .A3(_06387_),
    .A4(_06388_),
    .ZN(_06389_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13292_ (.I(_06389_),
    .Z(_06390_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13293_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[9] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ),
    .S(_03499_),
    .Z(_06391_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _13294_ (.A1(_06281_),
    .A2(_06284_),
    .A3(_06391_),
    .ZN(_06392_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13295_ (.I(_06392_),
    .ZN(_06393_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13296_ (.A1(_06313_),
    .A2(_06393_),
    .B(_06389_),
    .ZN(_06394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13297_ (.I(_06301_),
    .Z(_06395_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _13298_ (.A1(_06289_),
    .A2(_06390_),
    .B1(_06394_),
    .B2(_06373_),
    .C(_06395_),
    .ZN(_06396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13299_ (.I(_06328_),
    .Z(_06397_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13300_ (.I(_06397_),
    .Z(_06398_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _13301_ (.A1(_06383_),
    .A2(_06362_),
    .B1(_06375_),
    .B2(_06396_),
    .C(_06398_),
    .ZN(_06399_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _13302_ (.A1(_06366_),
    .A2(_06376_),
    .B(_06381_),
    .C(_06399_),
    .ZN(_06400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13303_ (.I(_06130_),
    .Z(_06401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13304_ (.A1(_06118_),
    .A2(_06300_),
    .ZN(_06402_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13305_ (.I(_06402_),
    .Z(_06403_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13306_ (.I(_06387_),
    .Z(_06404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13307_ (.A1(_06368_),
    .A2(_06404_),
    .ZN(_06405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13308_ (.A1(_06374_),
    .A2(_06362_),
    .ZN(_06406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13309_ (.A1(_06405_),
    .A2(_06406_),
    .ZN(_06407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13310_ (.A1(_06403_),
    .A2(_06407_),
    .ZN(_06408_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13311_ (.I(_06134_),
    .Z(_06409_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13312_ (.A1(_06401_),
    .A2(_06408_),
    .B(_06409_),
    .ZN(_06410_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13313_ (.A1(_06338_),
    .A2(_06363_),
    .B1(_06400_),
    .B2(_06410_),
    .ZN(_06411_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13314_ (.I(_06138_),
    .Z(_06412_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13315_ (.I(_06412_),
    .Z(_06413_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13316_ (.A1(\mod.u_cpu.cpu.immdec.imm11_7[1] ),
    .A2(_06413_),
    .B(_06357_),
    .ZN(_06414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13317_ (.A1(_03271_),
    .A2(_06358_),
    .B1(_06411_),
    .B2(_06414_),
    .ZN(_01206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13318_ (.I(_06138_),
    .Z(_06415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13319_ (.I(_06415_),
    .Z(_06416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13320_ (.I(_06313_),
    .Z(_06417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13321_ (.I(_06417_),
    .Z(_06418_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13322_ (.A1(_03664_),
    .A2(_06416_),
    .B1(_06339_),
    .B2(_06418_),
    .ZN(_06419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13323_ (.A1(\mod.u_cpu.cpu.immdec.imm11_7[1] ),
    .A2(_06358_),
    .ZN(_06420_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13324_ (.I(_06064_),
    .Z(_06421_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13325_ (.I(_06421_),
    .Z(_06422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13326_ (.I(_06130_),
    .Z(_06423_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13327_ (.I(_06385_),
    .Z(_06424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13328_ (.A1(_06298_),
    .A2(_06304_),
    .ZN(_06425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13329_ (.A1(_06425_),
    .A2(_06402_),
    .ZN(_06426_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13330_ (.A1(_06316_),
    .A2(_06426_),
    .ZN(_06427_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13331_ (.A1(_06424_),
    .A2(_06370_),
    .B1(_06427_),
    .B2(_06417_),
    .ZN(_06428_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13332_ (.A1(_06417_),
    .A2(_06326_),
    .B(_06330_),
    .ZN(_06429_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13333_ (.A1(_06318_),
    .A2(_06428_),
    .B(_06429_),
    .ZN(_06430_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13334_ (.I(_06133_),
    .Z(_06431_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13335_ (.I(_06431_),
    .Z(_06432_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13336_ (.A1(_06423_),
    .A2(_06430_),
    .B(_06432_),
    .ZN(_06433_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13337_ (.I(_06125_),
    .Z(_06434_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13338_ (.I(_06379_),
    .Z(_06435_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13339_ (.A1(_06434_),
    .A2(_06435_),
    .ZN(_06436_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13340_ (.I(_06436_),
    .Z(_06437_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13341_ (.I(_06374_),
    .Z(_06438_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13342_ (.A1(_06438_),
    .A2(_06390_),
    .ZN(_06439_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _13343_ (.A1(_06437_),
    .A2(_06418_),
    .A3(_06403_),
    .A4(_06439_),
    .ZN(_06440_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13344_ (.I(_06121_),
    .Z(_06441_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13345_ (.I(_06441_),
    .Z(_06442_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13346_ (.I(_06424_),
    .Z(_06443_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13347_ (.A1(_06442_),
    .A2(_06314_),
    .B1(_06443_),
    .B2(_06382_),
    .ZN(_06444_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13348_ (.A1(_06433_),
    .A2(_06440_),
    .B1(_06444_),
    .B2(_06401_),
    .ZN(_06445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13349_ (.A1(_06422_),
    .A2(_06445_),
    .ZN(_06446_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _13350_ (.A1(_06358_),
    .A2(_06419_),
    .B(_06420_),
    .C(_06446_),
    .ZN(_01207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13351_ (.A1(_06441_),
    .A2(_06390_),
    .ZN(_06447_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13352_ (.I(_06316_),
    .Z(_06448_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13353_ (.I(_06448_),
    .Z(_06449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13354_ (.A1(_06434_),
    .A2(_06435_),
    .ZN(_06450_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13355_ (.I(_06450_),
    .Z(_06451_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13356_ (.I(_06426_),
    .Z(_06452_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _13357_ (.A1(_06449_),
    .A2(_06451_),
    .A3(_06452_),
    .ZN(_06453_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13358_ (.A1(_06395_),
    .A2(_06380_),
    .B(_06131_),
    .ZN(_06454_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13359_ (.I(_06454_),
    .Z(_06455_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13360_ (.I(_06455_),
    .Z(_06456_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _13361_ (.A1(_06437_),
    .A2(_06447_),
    .B(_06453_),
    .C(_06456_),
    .ZN(_06457_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13362_ (.I(_06391_),
    .Z(_06458_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13363_ (.I(_06458_),
    .Z(_06459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13364_ (.A1(_06422_),
    .A2(_06459_),
    .ZN(_06460_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13365_ (.I0(_03664_),
    .I1(_03663_),
    .S(_06356_),
    .Z(_06461_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13366_ (.A1(_06326_),
    .A2(_06391_),
    .B(_06330_),
    .ZN(_06462_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13367_ (.I(_06308_),
    .Z(_06463_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13368_ (.I(_06388_),
    .Z(_06464_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13369_ (.I(_06464_),
    .Z(_06465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13370_ (.I(_06369_),
    .Z(_06466_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13371_ (.A1(_06463_),
    .A2(_06448_),
    .B1(_06465_),
    .B2(_06466_),
    .ZN(_06467_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13372_ (.I(_06292_),
    .Z(_06468_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13373_ (.A1(_06468_),
    .A2(_06403_),
    .ZN(_06469_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _13374_ (.I(_06374_),
    .Z(_06470_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13375_ (.I(_06470_),
    .Z(_06471_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13376_ (.I(_06130_),
    .Z(_06472_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _13377_ (.A1(_06471_),
    .A2(_06464_),
    .B1(_06458_),
    .B2(_06395_),
    .C(_06472_),
    .ZN(_06473_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _13378_ (.A1(_06462_),
    .A2(_06467_),
    .B1(_06469_),
    .B2(_06473_),
    .ZN(_06474_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13379_ (.I(_06454_),
    .Z(_06475_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13380_ (.A1(_06139_),
    .A2(_06475_),
    .ZN(_06476_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13381_ (.A1(_06413_),
    .A2(_06461_),
    .B1(_06474_),
    .B2(_06476_),
    .ZN(_06477_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13382_ (.A1(_06457_),
    .A2(_06460_),
    .B(_06477_),
    .ZN(_01208_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _13383_ (.A1(_03665_),
    .A2(_03391_),
    .A3(_03672_),
    .ZN(_06478_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13384_ (.A1(_03663_),
    .A2(_06356_),
    .B(_06416_),
    .ZN(_06479_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13385_ (.A1(_06397_),
    .A2(_06129_),
    .ZN(_06480_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13386_ (.A1(_06480_),
    .A2(_06447_),
    .ZN(_06481_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13387_ (.I(_06064_),
    .Z(_06482_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13388_ (.I(_06482_),
    .Z(_06483_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13389_ (.A1(_06377_),
    .A2(_03449_),
    .Z(_06484_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13390_ (.A1(_05784_),
    .A2(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[10] ),
    .B(_06484_),
    .ZN(_06485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13391_ (.I(_06435_),
    .Z(_06486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13392_ (.A1(_06470_),
    .A2(_06397_),
    .ZN(_06487_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _13393_ (.A1(_06442_),
    .A2(_06398_),
    .B(_06486_),
    .C(_06487_),
    .ZN(_06488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13394_ (.A1(_06485_),
    .A2(_06488_),
    .ZN(_06489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13395_ (.A1(_06310_),
    .A2(_06329_),
    .ZN(_06490_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13396_ (.A1(_06483_),
    .A2(_06489_),
    .A3(_06490_),
    .ZN(_06491_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _13397_ (.A1(_06478_),
    .A2(_06479_),
    .B1(_06481_),
    .B2(_06491_),
    .ZN(_01209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13398_ (.I(_06285_),
    .Z(_06492_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13399_ (.I(_06310_),
    .Z(_06493_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13400_ (.I(_06434_),
    .Z(_06494_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13401_ (.A1(_06438_),
    .A2(_06493_),
    .B(_06494_),
    .ZN(_06495_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13402_ (.A1(_06381_),
    .A2(_06439_),
    .A3(_06495_),
    .ZN(_06496_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13403_ (.A1(_06432_),
    .A2(_06403_),
    .A3(_06496_),
    .ZN(_06497_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13404_ (.A1(_06483_),
    .A2(_06492_),
    .A3(_06497_),
    .ZN(_06498_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13405_ (.A1(\mod.u_cpu.cpu.immdec.imm30_25[0] ),
    .A2(_06413_),
    .B(_06357_),
    .ZN(_06499_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13406_ (.A1(_04223_),
    .A2(_06358_),
    .B1(_06498_),
    .B2(_06499_),
    .ZN(_01210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13407_ (.A1(_03790_),
    .A2(_06344_),
    .ZN(_06500_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13408_ (.I0(_06351_),
    .I1(\mod.u_cpu.rf_ram.memory[91][0] ),
    .S(_06500_),
    .Z(_06501_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13409_ (.I(_06501_),
    .Z(_01211_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13410_ (.I0(_06354_),
    .I1(\mod.u_cpu.rf_ram.memory[91][1] ),
    .S(_06500_),
    .Z(_06502_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13411_ (.I(_06502_),
    .Z(_01212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13412_ (.A1(_03910_),
    .A2(_06011_),
    .ZN(_06503_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13413_ (.I0(_06351_),
    .I1(\mod.u_cpu.rf_ram.memory[139][0] ),
    .S(_06503_),
    .Z(_06504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13414_ (.I(_06504_),
    .Z(_01213_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13415_ (.I0(_06354_),
    .I1(\mod.u_cpu.rf_ram.memory[139][1] ),
    .S(_06503_),
    .Z(_06505_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13416_ (.I(_06505_),
    .Z(_01214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13417_ (.A1(_05732_),
    .A2(_04847_),
    .ZN(_06506_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13418_ (.I0(_06351_),
    .I1(\mod.u_cpu.rf_ram.memory[339][0] ),
    .S(_06506_),
    .Z(_06507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13419_ (.I(_06507_),
    .Z(_01215_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13420_ (.I0(_06354_),
    .I1(\mod.u_cpu.rf_ram.memory[339][1] ),
    .S(_06506_),
    .Z(_06508_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13421_ (.I(_06508_),
    .Z(_01216_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13422_ (.A1(_03377_),
    .A2(_03668_),
    .B(net5),
    .ZN(_06509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13423_ (.I(_06509_),
    .Z(_06510_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13424_ (.I(_06510_),
    .Z(_06511_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13425_ (.A1(net5),
    .A2(_03677_),
    .ZN(_06512_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13426_ (.I(_06512_),
    .Z(_06513_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13427_ (.I(_06513_),
    .Z(_06514_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13428_ (.A1(_03371_),
    .A2(_06511_),
    .B1(_06514_),
    .B2(_03492_),
    .ZN(_06515_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13429_ (.I(_06515_),
    .ZN(_01217_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13430_ (.A1(_03492_),
    .A2(_06511_),
    .B1(_06514_),
    .B2(_03508_),
    .ZN(_06516_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13431_ (.I(_06516_),
    .ZN(_01218_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13432_ (.A1(_03508_),
    .A2(_06511_),
    .B1(_06514_),
    .B2(_03507_),
    .ZN(_06517_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13433_ (.I(_06517_),
    .ZN(_01219_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13434_ (.A1(_03507_),
    .A2(_06511_),
    .B1(_06514_),
    .B2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[4] ),
    .ZN(_06518_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13435_ (.I(_06518_),
    .ZN(_01220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13436_ (.I(_06510_),
    .Z(_06519_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13437_ (.I(_06513_),
    .Z(_06520_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13438_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[4] ),
    .A2(_06519_),
    .B1(_06520_),
    .B2(_03520_),
    .ZN(_06521_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13439_ (.I(_06521_),
    .ZN(_01221_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13440_ (.A1(_03520_),
    .A2(_06519_),
    .B1(_06520_),
    .B2(_03524_),
    .ZN(_06522_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13441_ (.I(_06522_),
    .ZN(_01222_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13442_ (.A1(_03524_),
    .A2(_06519_),
    .B1(_06520_),
    .B2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[7] ),
    .ZN(_06523_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13443_ (.I(_06523_),
    .ZN(_01223_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13444_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[7] ),
    .A2(_06519_),
    .B1(_06520_),
    .B2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[8] ),
    .ZN(_06524_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13445_ (.I(_06524_),
    .ZN(_01224_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13446_ (.I(_06510_),
    .Z(_06525_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13447_ (.I(_06513_),
    .Z(_06526_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13448_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[8] ),
    .A2(_06525_),
    .B1(_06526_),
    .B2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[9] ),
    .ZN(_06527_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13449_ (.I(_06527_),
    .ZN(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13450_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[9] ),
    .A2(_06525_),
    .B1(_06526_),
    .B2(_03541_),
    .ZN(_06528_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13451_ (.I(_06528_),
    .ZN(_01226_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13452_ (.A1(_03541_),
    .A2(_06525_),
    .B1(_06526_),
    .B2(_03547_),
    .ZN(_06529_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13453_ (.I(_06529_),
    .ZN(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13454_ (.A1(_03547_),
    .A2(_06525_),
    .B1(_06526_),
    .B2(_03552_),
    .ZN(_06530_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13455_ (.I(_06530_),
    .ZN(_01228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13456_ (.I(_06510_),
    .Z(_06531_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13457_ (.I(_06513_),
    .Z(_06532_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13458_ (.A1(_03552_),
    .A2(_06531_),
    .B1(_06532_),
    .B2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[13] ),
    .ZN(_06533_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13459_ (.I(_06533_),
    .ZN(_01229_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13460_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[13] ),
    .A2(_06531_),
    .B1(_06532_),
    .B2(_03569_),
    .ZN(_06534_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13461_ (.I(_06534_),
    .ZN(_01230_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13462_ (.A1(_03569_),
    .A2(_06531_),
    .B1(_06532_),
    .B2(_03574_),
    .ZN(_06535_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13463_ (.I(_06535_),
    .ZN(_01231_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13464_ (.A1(_03574_),
    .A2(_06531_),
    .B1(_06532_),
    .B2(_03578_),
    .ZN(_06536_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13465_ (.I(_06536_),
    .ZN(_01232_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13466_ (.I(_06509_),
    .Z(_06537_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13467_ (.I(_06537_),
    .Z(_06538_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13468_ (.I(_06512_),
    .Z(_06539_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13469_ (.I(_06539_),
    .Z(_06540_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13470_ (.A1(_03578_),
    .A2(_06538_),
    .B1(_06540_),
    .B2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[17] ),
    .ZN(_06541_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13471_ (.I(_06541_),
    .ZN(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13472_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[17] ),
    .A2(_06538_),
    .B1(_06540_),
    .B2(_03588_),
    .ZN(_06542_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13473_ (.I(_06542_),
    .ZN(_01234_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13474_ (.A1(_03588_),
    .A2(_06538_),
    .B1(_06540_),
    .B2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[19] ),
    .ZN(_06543_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13475_ (.I(_06543_),
    .ZN(_01235_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13476_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[19] ),
    .A2(_06538_),
    .B1(_06540_),
    .B2(_03598_),
    .ZN(_06544_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13477_ (.I(_06544_),
    .ZN(_01236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13478_ (.I(_06537_),
    .Z(_06545_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13479_ (.I(_06539_),
    .Z(_06546_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13480_ (.A1(_03598_),
    .A2(_06545_),
    .B1(_06546_),
    .B2(_03602_),
    .ZN(_06547_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13481_ (.I(_06547_),
    .ZN(_01237_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13482_ (.A1(_03602_),
    .A2(_06545_),
    .B1(_06546_),
    .B2(_03605_),
    .ZN(_06548_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13483_ (.I(_06548_),
    .ZN(_01238_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13484_ (.A1(_03605_),
    .A2(_06545_),
    .B1(_06546_),
    .B2(_03610_),
    .ZN(_06549_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13485_ (.I(_06549_),
    .ZN(_01239_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13486_ (.A1(_03610_),
    .A2(_06545_),
    .B1(_06546_),
    .B2(_03616_),
    .ZN(_06550_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13487_ (.I(_06550_),
    .ZN(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13488_ (.I(_06537_),
    .Z(_06551_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13489_ (.I(_06539_),
    .Z(_06552_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13490_ (.A1(_03616_),
    .A2(_06551_),
    .B1(_06552_),
    .B2(_03624_),
    .ZN(_06553_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13491_ (.I(_06553_),
    .ZN(_01241_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13492_ (.A1(_03624_),
    .A2(_06551_),
    .B1(_06552_),
    .B2(_03631_),
    .ZN(_06554_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13493_ (.I(_06554_),
    .ZN(_01242_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13494_ (.A1(_03631_),
    .A2(_06551_),
    .B1(_06552_),
    .B2(_03635_),
    .ZN(_06555_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13495_ (.I(_06555_),
    .ZN(_01243_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13496_ (.A1(_03635_),
    .A2(_06551_),
    .B1(_06552_),
    .B2(_03642_),
    .ZN(_06556_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13497_ (.I(_06556_),
    .ZN(_01244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13498_ (.I(_06537_),
    .Z(_06557_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13499_ (.I(_06539_),
    .Z(_06558_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13500_ (.A1(_03642_),
    .A2(_06557_),
    .B1(_06558_),
    .B2(_03648_),
    .ZN(_06559_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13501_ (.I(_06559_),
    .ZN(_01245_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13502_ (.A1(_03648_),
    .A2(_06557_),
    .B1(_06558_),
    .B2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[30] ),
    .ZN(_06560_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13503_ (.I(_06560_),
    .ZN(_01246_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13504_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[30] ),
    .A2(_06557_),
    .B1(_06558_),
    .B2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[31] ),
    .ZN(_06561_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13505_ (.I(_06561_),
    .ZN(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13506_ (.A1(_06142_),
    .A2(_03250_),
    .ZN(_06562_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13507_ (.A1(\mod.u_cpu.cpu.ctrl.i_jump ),
    .A2(_03296_),
    .B(_06562_),
    .ZN(_06563_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13508_ (.A1(\mod.u_cpu.cpu.ctrl.i_jump ),
    .A2(_03325_),
    .B(_06563_),
    .ZN(_06564_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13509_ (.A1(_06562_),
    .A2(_03302_),
    .A3(_03260_),
    .ZN(_06565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13510_ (.A1(_06564_),
    .A2(_06565_),
    .ZN(_06566_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13511_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[31] ),
    .A2(_06557_),
    .B1(_06558_),
    .B2(_06566_),
    .ZN(_06567_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13512_ (.I(_06567_),
    .ZN(_01248_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13513_ (.I(_05791_),
    .Z(_06568_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _13514_ (.A1(\mod.u_cpu.cpu.state.o_cnt_r[1] ),
    .A2(_03388_),
    .B(_03337_),
    .C(_06568_),
    .ZN(_06569_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _13515_ (.A1(_03693_),
    .A2(_06568_),
    .B(_06569_),
    .ZN(_06570_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13516_ (.A1(_03426_),
    .A2(_06570_),
    .ZN(_06571_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13517_ (.A1(_03425_),
    .A2(_06570_),
    .B(_06571_),
    .ZN(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13518_ (.A1(_03685_),
    .A2(_03690_),
    .Z(_06572_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13519_ (.A1(_06568_),
    .A2(_03691_),
    .A3(_06572_),
    .ZN(_06573_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13520_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_adr[2] ),
    .A2(_03669_),
    .ZN(_06574_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13521_ (.A1(_06573_),
    .A2(_06574_),
    .ZN(_06575_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13522_ (.I0(_03426_),
    .I1(_06575_),
    .S(_06570_),
    .Z(_06576_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13523_ (.I(_06576_),
    .Z(_01250_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13524_ (.I(_03923_),
    .Z(_06577_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13525_ (.I(_06577_),
    .Z(_06578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13526_ (.A1(_03980_),
    .A2(_05373_),
    .ZN(_06579_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13527_ (.I0(_06578_),
    .I1(\mod.u_cpu.rf_ram.memory[129][0] ),
    .S(_06579_),
    .Z(_06580_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13528_ (.I(_06580_),
    .Z(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13529_ (.I(_06236_),
    .Z(_06581_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13530_ (.I0(_06581_),
    .I1(\mod.u_cpu.rf_ram.memory[129][1] ),
    .S(_06579_),
    .Z(_06582_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13531_ (.I(_06582_),
    .Z(_01252_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13532_ (.I(_03292_),
    .Z(_06583_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13533_ (.I(_06583_),
    .Z(_06584_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13534_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[2] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[3] ),
    .S(_06584_),
    .Z(_06585_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13535_ (.I(_06585_),
    .Z(_01253_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13536_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[3] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[4] ),
    .S(_06584_),
    .Z(_06586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13537_ (.I(_06586_),
    .Z(_01254_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13538_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[4] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[5] ),
    .S(_06584_),
    .Z(_06587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13539_ (.I(_06587_),
    .Z(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13540_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[5] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[6] ),
    .S(_06584_),
    .Z(_06588_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13541_ (.I(_06588_),
    .Z(_01256_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13542_ (.I(_06583_),
    .Z(_06589_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13543_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[6] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[7] ),
    .S(_06589_),
    .Z(_06590_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13544_ (.I(_06590_),
    .Z(_01257_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13545_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[7] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[8] ),
    .S(_06589_),
    .Z(_06591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13546_ (.I(_06591_),
    .Z(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13547_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[8] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[9] ),
    .S(_06589_),
    .Z(_06592_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13548_ (.I(_06592_),
    .Z(_01259_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13549_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[9] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[10] ),
    .S(_06589_),
    .Z(_06593_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13550_ (.I(_06593_),
    .Z(_01260_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13551_ (.I(_06583_),
    .Z(_06594_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13552_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[10] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[11] ),
    .S(_06594_),
    .Z(_06595_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13553_ (.I(_06595_),
    .Z(_01261_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13554_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[11] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[12] ),
    .S(_06594_),
    .Z(_06596_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13555_ (.I(_06596_),
    .Z(_01262_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13556_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[12] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[13] ),
    .S(_06594_),
    .Z(_06597_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13557_ (.I(_06597_),
    .Z(_01263_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13558_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[13] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[14] ),
    .S(_06594_),
    .Z(_06598_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13559_ (.I(_06598_),
    .Z(_01264_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13560_ (.I(_06583_),
    .Z(_06599_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13561_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[14] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[15] ),
    .S(_06599_),
    .Z(_06600_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13562_ (.I(_06600_),
    .Z(_01265_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13563_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[15] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[16] ),
    .S(_06599_),
    .Z(_06601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13564_ (.I(_06601_),
    .Z(_01266_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13565_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[16] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[17] ),
    .S(_06599_),
    .Z(_06602_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13566_ (.I(_06602_),
    .Z(_01267_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13567_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[17] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[18] ),
    .S(_06599_),
    .Z(_06603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13568_ (.I(_06603_),
    .Z(_01268_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13569_ (.I(_03692_),
    .Z(_06604_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13570_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[18] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[19] ),
    .S(_06604_),
    .Z(_06605_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13571_ (.I(_06605_),
    .Z(_01269_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13572_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[19] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[20] ),
    .S(_06604_),
    .Z(_06606_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13573_ (.I(_06606_),
    .Z(_01270_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13574_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[20] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[21] ),
    .S(_06604_),
    .Z(_06607_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13575_ (.I(_06607_),
    .Z(_01271_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13576_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[21] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[22] ),
    .S(_06604_),
    .Z(_06608_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13577_ (.I(_06608_),
    .Z(_01272_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13578_ (.I(_03692_),
    .Z(_06609_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13579_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[22] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[23] ),
    .S(_06609_),
    .Z(_06610_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13580_ (.I(_06610_),
    .Z(_01273_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13581_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[23] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[24] ),
    .S(_06609_),
    .Z(_06611_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13582_ (.I(_06611_),
    .Z(_01274_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13583_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[24] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[25] ),
    .S(_06609_),
    .Z(_06612_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13584_ (.I(_06612_),
    .Z(_01275_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13585_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[25] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[26] ),
    .S(_06609_),
    .Z(_06613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13586_ (.I(_06613_),
    .Z(_01276_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13587_ (.I(_03692_),
    .Z(_06614_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13588_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[26] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[27] ),
    .S(_06614_),
    .Z(_06615_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13589_ (.I(_06615_),
    .Z(_01277_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13590_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[27] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[28] ),
    .S(_06614_),
    .Z(_06616_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13591_ (.I(_06616_),
    .Z(_01278_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13592_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[28] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[29] ),
    .S(_06614_),
    .Z(_06617_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13593_ (.I(_06617_),
    .Z(_01279_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13594_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[29] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[30] ),
    .S(_06614_),
    .Z(_06618_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13595_ (.I(_06618_),
    .Z(_01280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13596_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_adr[30] ),
    .A2(_03694_),
    .ZN(_06619_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13597_ (.A1(_03659_),
    .A2(_03694_),
    .B(_06619_),
    .ZN(_01281_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13598_ (.A1(\mod.u_cpu.cpu.bufreg.i_sh_signed ),
    .A2(_03669_),
    .B(_03693_),
    .ZN(_06620_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _13599_ (.A1(_03694_),
    .A2(_06573_),
    .B1(_06620_),
    .B2(_03659_),
    .ZN(_01282_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _13600_ (.A1(_03713_),
    .A2(_04922_),
    .ZN(_06621_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13601_ (.I0(\mod.u_cpu.rf_ram.memory[329][0] ),
    .I1(_03899_),
    .S(_06621_),
    .Z(_06622_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13602_ (.I(_06622_),
    .Z(_01283_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13603_ (.I0(\mod.u_cpu.rf_ram.memory[329][1] ),
    .I1(_06221_),
    .S(_06621_),
    .Z(_06623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13604_ (.I(_06623_),
    .Z(_01284_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13605_ (.A1(_03362_),
    .A2(_03354_),
    .ZN(_06624_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13606_ (.A1(_01429_),
    .A2(_03307_),
    .B(_03315_),
    .ZN(_06625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13607_ (.A1(_03309_),
    .A2(_06625_),
    .ZN(_06626_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13608_ (.A1(_03381_),
    .A2(_06626_),
    .Z(_06627_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13609_ (.A1(_03365_),
    .A2(_06625_),
    .B(_06627_),
    .ZN(_06628_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _13610_ (.A1(_03365_),
    .A2(_06625_),
    .A3(_06627_),
    .Z(_06629_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _13611_ (.A1(\mod.u_cpu.cpu.alu.cmp_r ),
    .A2(_03687_),
    .B(_03305_),
    .C(_06624_),
    .ZN(_06630_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _13612_ (.A1(_06624_),
    .A2(_06628_),
    .A3(_06629_),
    .B(_06630_),
    .ZN(_06631_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13613_ (.A1(_03378_),
    .A2(_06631_),
    .ZN(_06632_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13614_ (.A1(_03313_),
    .A2(_03378_),
    .B(_06632_),
    .ZN(_01285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13615_ (.A1(_04844_),
    .A2(_05020_),
    .ZN(_06633_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13616_ (.A1(_06249_),
    .A2(_06633_),
    .ZN(_06634_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13617_ (.A1(_01926_),
    .A2(_06633_),
    .B(_06634_),
    .ZN(_01286_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13618_ (.I0(_06581_),
    .I1(\mod.u_cpu.rf_ram.memory[319][1] ),
    .S(_06633_),
    .Z(_06635_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13619_ (.I(_06635_),
    .Z(_01287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13620_ (.A1(_05164_),
    .A2(_04989_),
    .ZN(_06636_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13621_ (.A1(_06249_),
    .A2(_06636_),
    .ZN(_06637_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13622_ (.A1(_01935_),
    .A2(_06636_),
    .B(_06637_),
    .ZN(_01288_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13623_ (.I0(_06581_),
    .I1(\mod.u_cpu.rf_ram.memory[309][1] ),
    .S(_06636_),
    .Z(_06638_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13624_ (.I(_06638_),
    .Z(_01289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13625_ (.A1(\mod.u_cpu.cpu.genblk3.csr.timer_irq_r ),
    .A2(_06111_),
    .ZN(_06639_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13626_ (.A1(_06111_),
    .A2(_06112_),
    .B(_06639_),
    .ZN(_01290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13627_ (.I(_06415_),
    .Z(_06640_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13628_ (.I(_06640_),
    .Z(_06641_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13629_ (.I(_06332_),
    .ZN(_06642_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _13630_ (.A1(_06485_),
    .A2(_06284_),
    .A3(_06322_),
    .A4(_06305_),
    .ZN(_06643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13631_ (.A1(_06371_),
    .A2(_06310_),
    .ZN(_06644_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _13632_ (.A1(_06319_),
    .A2(_06324_),
    .A3(_06643_),
    .A4(_06644_),
    .ZN(_06645_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13633_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[31] ),
    .I1(_03458_),
    .S(_03503_),
    .Z(_06646_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13634_ (.I(_06455_),
    .Z(_06647_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13635_ (.A1(_06642_),
    .A2(_06645_),
    .B1(_06646_),
    .B2(_06647_),
    .ZN(_06648_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13636_ (.I(_06412_),
    .Z(_06649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13637_ (.A1(\mod.u_cpu.cpu.immdec.imm31 ),
    .A2(_06649_),
    .ZN(_06650_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13638_ (.A1(_06641_),
    .A2(_06648_),
    .B(_06650_),
    .ZN(_01291_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13639_ (.I(\mod.u_cpu.cpu.immdec.imm19_12_20[0] ),
    .ZN(_06651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13640_ (.A1(_03297_),
    .A2(_03681_),
    .ZN(_06652_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13641_ (.A1(_03297_),
    .A2(\mod.u_cpu.cpu.decode.opcode[1] ),
    .B(_06652_),
    .ZN(_06653_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13642_ (.A1(_03274_),
    .A2(_06653_),
    .Z(_06654_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13643_ (.A1(_03390_),
    .A2(_06654_),
    .B(_06137_),
    .ZN(_06655_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13644_ (.I(_06655_),
    .Z(_06656_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13645_ (.I(_06656_),
    .Z(_06657_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13646_ (.I(_06655_),
    .Z(_06658_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13647_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[20] ),
    .I1(\mod.u_arbiter.i_wb_cpu_rdt[4] ),
    .S(_06334_),
    .Z(_06659_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _13648_ (.A1(_06289_),
    .A2(_06313_),
    .A3(_06361_),
    .A4(_06393_),
    .Z(_06660_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13649_ (.I(_06404_),
    .Z(_06661_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13650_ (.A1(_06320_),
    .A2(_06368_),
    .ZN(_06662_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13651_ (.A1(_06661_),
    .A2(_06662_),
    .ZN(_06663_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13652_ (.I(_06129_),
    .Z(_06664_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _13653_ (.A1(_06447_),
    .A2(_06660_),
    .B(_06663_),
    .C(_06664_),
    .ZN(_06665_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13654_ (.A1(_06298_),
    .A2(_06299_),
    .ZN(_06666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13655_ (.A1(_06304_),
    .A2(_06666_),
    .ZN(_06667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13656_ (.A1(_06312_),
    .A2(_06392_),
    .ZN(_06668_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13657_ (.A1(_06361_),
    .A2(_06668_),
    .ZN(_06669_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13658_ (.A1(_06667_),
    .A2(_06669_),
    .ZN(_06670_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13659_ (.A1(_06371_),
    .A2(_06670_),
    .ZN(_06671_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13660_ (.I(_06671_),
    .Z(_06672_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13661_ (.A1(_06309_),
    .A2(_06404_),
    .A3(_06402_),
    .ZN(_06673_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _13662_ (.A1(_06434_),
    .A2(_06644_),
    .A3(_06673_),
    .Z(_06674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13663_ (.A1(_06661_),
    .A2(_06369_),
    .ZN(_06675_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _13664_ (.A1(_06672_),
    .A2(_06674_),
    .B1(_06675_),
    .B2(_06472_),
    .C(_06134_),
    .ZN(_06676_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _13665_ (.A1(_06338_),
    .A2(_06659_),
    .B1(_06665_),
    .B2(_06676_),
    .ZN(_06677_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13666_ (.I(_06415_),
    .Z(_06678_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13667_ (.A1(\mod.u_cpu.cpu.immdec.imm19_12_20[1] ),
    .A2(_06678_),
    .ZN(_06679_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13668_ (.A1(_06677_),
    .A2(_06679_),
    .ZN(_06680_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13669_ (.A1(_06658_),
    .A2(_06680_),
    .ZN(_06681_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13670_ (.A1(_06651_),
    .A2(_06657_),
    .B(_06681_),
    .ZN(_01292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13671_ (.I(_06670_),
    .Z(_06682_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13672_ (.I(_06291_),
    .Z(_06683_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _13673_ (.A1(_06683_),
    .A2(_06293_),
    .B(_06282_),
    .C(_06294_),
    .ZN(_06684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _13674_ (.A1(_06304_),
    .A2(_06370_),
    .B1(_06682_),
    .B2(_06661_),
    .C1(_06684_),
    .C2(_06306_),
    .ZN(_06685_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13675_ (.A1(_06431_),
    .A2(_06490_),
    .ZN(_06686_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13676_ (.A1(_06437_),
    .A2(_06448_),
    .B1(_06686_),
    .B2(_06372_),
    .ZN(_06687_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13677_ (.A1(_06451_),
    .A2(_06685_),
    .B(_06687_),
    .ZN(_06688_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13678_ (.A1(_06421_),
    .A2(_06688_),
    .ZN(_06689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13679_ (.A1(\mod.u_cpu.cpu.immdec.imm19_12_20[2] ),
    .A2(_06678_),
    .ZN(_06690_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13680_ (.A1(_06689_),
    .A2(_06690_),
    .ZN(_06691_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13681_ (.I0(\mod.u_cpu.cpu.immdec.imm19_12_20[1] ),
    .I1(_06691_),
    .S(_06658_),
    .Z(_06692_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13682_ (.I(_06692_),
    .Z(_01293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13683_ (.A1(_06482_),
    .A2(_06475_),
    .ZN(_06693_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13684_ (.I(_06367_),
    .Z(_06694_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13685_ (.A1(_06694_),
    .A2(_06398_),
    .ZN(_06695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13686_ (.A1(_06424_),
    .A2(_06682_),
    .ZN(_06696_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _13687_ (.A1(_06292_),
    .A2(_06485_),
    .B(_06294_),
    .C(_06305_),
    .ZN(_06697_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _13688_ (.A1(_06494_),
    .A2(_06644_),
    .A3(_06696_),
    .A4(_06697_),
    .ZN(_06698_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13689_ (.A1(_06695_),
    .A2(_06698_),
    .ZN(_06699_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _13690_ (.A1(_06693_),
    .A2(_06463_),
    .B1(_06699_),
    .B2(_06409_),
    .ZN(_06700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13691_ (.A1(\mod.u_cpu.cpu.immdec.imm19_12_20[3] ),
    .A2(_06678_),
    .ZN(_06701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13692_ (.A1(_06656_),
    .A2(_06701_),
    .ZN(_06702_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _13693_ (.A1(\mod.u_cpu.cpu.immdec.imm19_12_20[2] ),
    .A2(_06658_),
    .B1(_06700_),
    .B2(_06702_),
    .ZN(_06703_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13694_ (.I(_06703_),
    .ZN(_01294_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13695_ (.I(_05787_),
    .Z(_06704_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _13696_ (.A1(_06295_),
    .A2(_06306_),
    .B1(_06464_),
    .B2(_06682_),
    .C1(_06493_),
    .C2(_06323_),
    .ZN(_06705_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _13697_ (.A1(_06694_),
    .A2(_06431_),
    .B1(_06450_),
    .B2(_06705_),
    .ZN(_06706_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13698_ (.A1(_06421_),
    .A2(_06706_),
    .ZN(_06707_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13699_ (.A1(_03364_),
    .A2(_06704_),
    .B(_06707_),
    .ZN(_06708_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13700_ (.I(_06655_),
    .Z(_06709_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13701_ (.I0(\mod.u_cpu.cpu.immdec.imm19_12_20[3] ),
    .I1(_06708_),
    .S(_06709_),
    .Z(_06710_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13702_ (.I(_06710_),
    .Z(_01295_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _13703_ (.A1(_06371_),
    .A2(_06389_),
    .ZN(_06711_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _13704_ (.A1(_06470_),
    .A2(_06711_),
    .B(_06480_),
    .C(_06320_),
    .ZN(_06712_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13705_ (.A1(_06317_),
    .A2(_06644_),
    .ZN(_06713_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13706_ (.I(_06669_),
    .Z(_06714_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _13707_ (.A1(_06683_),
    .A2(_06667_),
    .A3(_06714_),
    .B1(_06493_),
    .B2(_06406_),
    .ZN(_06715_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _13708_ (.A1(_06318_),
    .A2(_06364_),
    .B1(_06713_),
    .B2(_06715_),
    .C(_06365_),
    .ZN(_06716_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13709_ (.A1(_06380_),
    .A2(_06448_),
    .ZN(_06717_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13710_ (.A1(_06694_),
    .A2(_06363_),
    .B(_06717_),
    .ZN(_06718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13711_ (.A1(_06716_),
    .A2(_06718_),
    .ZN(_06719_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _13712_ (.A1(_06363_),
    .A2(_06712_),
    .B(_06719_),
    .C(_06135_),
    .ZN(_06720_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _13713_ (.A1(\mod.u_cpu.cpu.immdec.imm19_12_20[5] ),
    .A2(_06704_),
    .B1(_06471_),
    .B2(_06693_),
    .C(_06656_),
    .ZN(_06721_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _13714_ (.A1(_03364_),
    .A2(_06657_),
    .B1(_06720_),
    .B2(_06721_),
    .ZN(_01296_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13715_ (.I(\mod.u_cpu.cpu.immdec.imm19_12_20[5] ),
    .ZN(_06722_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13716_ (.I(_05784_),
    .Z(_06723_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13717_ (.A1(_06723_),
    .A2(\mod.u_arbiter.i_wb_cpu_rdt[16] ),
    .ZN(_06724_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13718_ (.A1(_06723_),
    .A2(_06123_),
    .B(_06724_),
    .ZN(_06725_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13719_ (.I(_06320_),
    .Z(_06726_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13720_ (.A1(_06726_),
    .A2(_06314_),
    .B1(_06725_),
    .B2(_06441_),
    .ZN(_06727_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13721_ (.A1(_06717_),
    .A2(_06727_),
    .B(_06475_),
    .ZN(_06728_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13722_ (.A1(_06463_),
    .A2(_06662_),
    .ZN(_06729_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13723_ (.A1(_06362_),
    .A2(_06668_),
    .B(_06293_),
    .ZN(_06730_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13724_ (.A1(_06382_),
    .A2(_06493_),
    .ZN(_06731_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _13725_ (.A1(_06729_),
    .A2(_06730_),
    .B1(_06731_),
    .B2(_06314_),
    .C(_06713_),
    .ZN(_06732_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13726_ (.A1(_06438_),
    .A2(_06711_),
    .ZN(_06733_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _13727_ (.A1(_06417_),
    .A2(_06733_),
    .B(_06321_),
    .C(_06486_),
    .ZN(_06734_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13728_ (.I(_06494_),
    .Z(_06735_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _13729_ (.A1(_06429_),
    .A2(_06732_),
    .B1(_06734_),
    .B2(_06735_),
    .ZN(_06736_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _13730_ (.A1(_06456_),
    .A2(_06725_),
    .B1(_06728_),
    .B2(_06736_),
    .C(_06640_),
    .ZN(_06737_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13731_ (.A1(\mod.u_cpu.cpu.immdec.imm19_12_20[6] ),
    .A2(_06483_),
    .B(_06709_),
    .ZN(_06738_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _13732_ (.A1(_06722_),
    .A2(_06657_),
    .B1(_06737_),
    .B2(_06738_),
    .ZN(_01297_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13733_ (.I(_06723_),
    .Z(_06739_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13734_ (.A1(_06723_),
    .A2(\mod.u_arbiter.i_wb_cpu_rdt[17] ),
    .ZN(_06740_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13735_ (.A1(_06739_),
    .A2(_03424_),
    .B(_06740_),
    .ZN(_06741_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _13736_ (.A1(_06726_),
    .A2(_06459_),
    .B1(_06741_),
    .B2(_06442_),
    .C(_06381_),
    .ZN(_06742_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _13737_ (.A1(_06288_),
    .A2(_06667_),
    .A3(_06669_),
    .ZN(_06743_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13738_ (.I(_06743_),
    .Z(_06744_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13739_ (.A1(_06713_),
    .A2(_06744_),
    .ZN(_06745_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13740_ (.A1(_06470_),
    .A2(_06425_),
    .A3(_06458_),
    .ZN(_06746_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13741_ (.A1(_06745_),
    .A2(_06746_),
    .B(_06462_),
    .ZN(_06747_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _13742_ (.A1(_06459_),
    .A2(_06712_),
    .B(_06747_),
    .C(_06423_),
    .ZN(_06748_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _13743_ (.A1(_06678_),
    .A2(_06456_),
    .A3(_06742_),
    .A4(_06748_),
    .ZN(_06749_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13744_ (.A1(\mod.u_cpu.cpu.immdec.imm19_12_20[7] ),
    .A2(_06139_),
    .B1(_06338_),
    .B2(_06741_),
    .ZN(_06750_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13745_ (.A1(_06656_),
    .A2(_06750_),
    .ZN(_06751_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _13746_ (.A1(\mod.u_cpu.cpu.immdec.imm19_12_20[6] ),
    .A2(_06658_),
    .B1(_06749_),
    .B2(_06751_),
    .ZN(_06752_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13747_ (.I(_06752_),
    .ZN(_01298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13748_ (.I(_06482_),
    .Z(_06753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13749_ (.A1(_06335_),
    .A2(_03428_),
    .ZN(_06754_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13750_ (.A1(_03510_),
    .A2(\mod.u_arbiter.i_wb_cpu_rdt[18] ),
    .B(_06754_),
    .ZN(_06755_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _13751_ (.A1(_06323_),
    .A2(_06425_),
    .B1(_06326_),
    .B2(_06281_),
    .C(_06330_),
    .ZN(_06756_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13752_ (.A1(_06666_),
    .A2(_06671_),
    .B(_06756_),
    .ZN(_06757_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _13753_ (.A1(_06726_),
    .A2(_06472_),
    .B1(_06283_),
    .B2(_06712_),
    .C(_06757_),
    .ZN(_06758_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _13754_ (.A1(_06432_),
    .A2(_06755_),
    .B(_06758_),
    .C(_06065_),
    .ZN(_06759_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _13755_ (.A1(\mod.u_cpu.cpu.immdec.imm19_12_20[8] ),
    .A2(_06753_),
    .B(_06709_),
    .C(_06759_),
    .ZN(_06760_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13756_ (.A1(_01479_),
    .A2(_06657_),
    .B(_06760_),
    .ZN(_01299_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _13757_ (.A1(_06492_),
    .A2(_06319_),
    .B1(_06713_),
    .B2(_06744_),
    .C(_06365_),
    .ZN(_06761_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13758_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[19] ),
    .I1(\mod.u_arbiter.i_wb_cpu_rdt[3] ),
    .S(_03509_),
    .Z(_06762_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _13759_ (.A1(_06492_),
    .A2(_06712_),
    .B1(_06762_),
    .B2(_06475_),
    .C(_06412_),
    .ZN(_06763_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13760_ (.A1(\mod.u_cpu.cpu.immdec.imm31 ),
    .A2(_03274_),
    .Z(_06764_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13761_ (.A1(_03686_),
    .A2(_06764_),
    .ZN(_06765_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13762_ (.A1(_03298_),
    .A2(\mod.u_cpu.cpu.immdec.imm24_20[0] ),
    .B(_06421_),
    .ZN(_06766_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13763_ (.A1(_06761_),
    .A2(_06763_),
    .B1(_06765_),
    .B2(_06766_),
    .ZN(_06767_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13764_ (.I0(\mod.u_cpu.cpu.immdec.imm19_12_20[8] ),
    .I1(_06767_),
    .S(_06709_),
    .Z(_06768_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13765_ (.I(_06768_),
    .Z(_01300_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13766_ (.A1(\mod.u_cpu.cpu.immdec.imm7 ),
    .A2(_06753_),
    .ZN(_06769_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13767_ (.A1(_06764_),
    .A2(_03391_),
    .B(_06416_),
    .ZN(_06770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13768_ (.A1(_03674_),
    .A2(_06769_),
    .B1(_06770_),
    .B2(_06411_),
    .ZN(_01301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13769_ (.A1(_03670_),
    .A2(_03396_),
    .ZN(_06771_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13770_ (.A1(_03403_),
    .A2(_06771_),
    .B(_03377_),
    .ZN(_06772_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13771_ (.A1(_06415_),
    .A2(_06772_),
    .Z(_06773_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13772_ (.I(_06773_),
    .Z(_06774_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13773_ (.A1(_06309_),
    .A2(_06666_),
    .ZN(_06775_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _13774_ (.A1(_06289_),
    .A2(_06775_),
    .B(_06643_),
    .C(_06317_),
    .ZN(_06776_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13775_ (.I(_06776_),
    .ZN(_06777_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13776_ (.A1(_06322_),
    .A2(_06714_),
    .ZN(_06778_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13777_ (.A1(_06667_),
    .A2(_06778_),
    .ZN(_06779_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _13778_ (.A1(_06404_),
    .A2(_06744_),
    .B1(_06779_),
    .B2(_06426_),
    .ZN(_06780_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13779_ (.A1(_06777_),
    .A2(_06780_),
    .B(_06331_),
    .ZN(_06781_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13780_ (.A1(_06494_),
    .A2(_06324_),
    .B(_06380_),
    .ZN(_06782_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _13781_ (.A1(_06381_),
    .A2(_06372_),
    .B1(_06781_),
    .B2(_06782_),
    .C(_06432_),
    .ZN(_06783_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13782_ (.A1(_03509_),
    .A2(\mod.u_arbiter.i_wb_cpu_rdt[25] ),
    .Z(_06784_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _13783_ (.A1(_06739_),
    .A2(\mod.u_arbiter.i_wb_cpu_rdt[9] ),
    .B(_06455_),
    .C(_06784_),
    .ZN(_06785_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13784_ (.A1(_06065_),
    .A2(_06783_),
    .A3(_06785_),
    .ZN(_06786_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13785_ (.A1(\mod.u_cpu.cpu.immdec.imm30_25[1] ),
    .A2(_06753_),
    .B(_06786_),
    .ZN(_06787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13786_ (.A1(\mod.u_cpu.cpu.immdec.imm30_25[0] ),
    .A2(_06774_),
    .ZN(_06788_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13787_ (.A1(_06774_),
    .A2(_06787_),
    .B(_06788_),
    .ZN(_01302_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13788_ (.I(\mod.u_cpu.cpu.immdec.imm30_25[1] ),
    .ZN(_06789_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13789_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[26] ),
    .I1(_03449_),
    .S(_03502_),
    .Z(_06790_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13790_ (.I(_06291_),
    .Z(_06791_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13791_ (.A1(_06791_),
    .A2(_06714_),
    .ZN(_06792_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _13792_ (.A1(_06425_),
    .A2(_06373_),
    .B1(_06402_),
    .B2(_06683_),
    .ZN(_06793_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _13793_ (.A1(_06779_),
    .A2(_06792_),
    .B(_06793_),
    .C(_06776_),
    .ZN(_06794_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13794_ (.A1(_06726_),
    .A2(_06407_),
    .B(_06486_),
    .ZN(_06795_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _13795_ (.A1(_06331_),
    .A2(_06794_),
    .B1(_06795_),
    .B2(_06735_),
    .ZN(_06796_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13796_ (.A1(_06321_),
    .A2(_06683_),
    .ZN(_06797_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _13797_ (.A1(_06383_),
    .A2(_06364_),
    .B1(_06790_),
    .B2(_06395_),
    .C(_06797_),
    .ZN(_06798_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13798_ (.A1(_06401_),
    .A2(_06798_),
    .B(_06409_),
    .ZN(_06799_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13799_ (.A1(_06339_),
    .A2(_06790_),
    .B1(_06796_),
    .B2(_06799_),
    .ZN(_06800_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13800_ (.A1(\mod.u_cpu.cpu.immdec.imm30_25[2] ),
    .A2(_06772_),
    .B(_06416_),
    .ZN(_06801_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13801_ (.A1(_06789_),
    .A2(_06774_),
    .B1(_06800_),
    .B2(_06801_),
    .ZN(_01303_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _13802_ (.A1(_06418_),
    .A2(_06466_),
    .B1(_06666_),
    .B2(_06443_),
    .C(_06486_),
    .ZN(_06802_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13803_ (.I(_06424_),
    .ZN(_06803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13804_ (.A1(_06803_),
    .A2(_06714_),
    .ZN(_06804_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _13805_ (.A1(_06468_),
    .A2(_06452_),
    .B1(_06779_),
    .B2(_06804_),
    .C(_06776_),
    .ZN(_06805_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _13806_ (.A1(_06735_),
    .A2(_06802_),
    .B1(_06805_),
    .B2(_06332_),
    .ZN(_06806_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13807_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[27] ),
    .I1(\mod.u_arbiter.i_wb_cpu_rdt[11] ),
    .S(_03509_),
    .Z(_06807_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13808_ (.A1(_06418_),
    .A2(_06449_),
    .B1(_06807_),
    .B2(_06442_),
    .ZN(_06808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13809_ (.A1(_06401_),
    .A2(_06808_),
    .ZN(_06809_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13810_ (.A1(_06476_),
    .A2(_06806_),
    .A3(_06809_),
    .ZN(_06810_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13811_ (.I(_06337_),
    .Z(_06811_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13812_ (.A1(_06482_),
    .A2(_06772_),
    .ZN(_06812_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _13813_ (.A1(\mod.u_cpu.cpu.immdec.imm30_25[2] ),
    .A2(_06773_),
    .B1(_06807_),
    .B2(_06811_),
    .C1(_06812_),
    .C2(\mod.u_cpu.cpu.immdec.imm30_25[3] ),
    .ZN(_06813_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13814_ (.A1(_06810_),
    .A2(_06813_),
    .ZN(_01304_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13815_ (.I(_06431_),
    .Z(_06814_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13816_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[28] ),
    .I1(\mod.u_arbiter.i_wb_cpu_rdt[12] ),
    .S(_03510_),
    .Z(_06815_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13817_ (.A1(_06423_),
    .A2(_06449_),
    .A3(_06459_),
    .ZN(_06816_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13818_ (.A1(_06814_),
    .A2(_06816_),
    .ZN(_06817_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _13819_ (.A1(_06363_),
    .A2(_06465_),
    .A3(_06668_),
    .B(_06779_),
    .ZN(_06818_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _13820_ (.A1(_06311_),
    .A2(_06458_),
    .B1(_06466_),
    .B2(_06372_),
    .C(_06776_),
    .ZN(_06819_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13821_ (.A1(_06818_),
    .A2(_06819_),
    .B(_06332_),
    .ZN(_06820_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _13822_ (.A1(_06814_),
    .A2(_06815_),
    .B1(_06817_),
    .B2(_06820_),
    .C(_06753_),
    .ZN(_06821_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13823_ (.A1(\mod.u_cpu.cpu.immdec.imm30_25[3] ),
    .A2(_06773_),
    .B1(_06812_),
    .B2(\mod.u_cpu.cpu.immdec.imm30_25[4] ),
    .ZN(_06822_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13824_ (.A1(_06821_),
    .A2(_06822_),
    .ZN(_01305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13825_ (.I(_06664_),
    .Z(_06823_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _13826_ (.A1(_06471_),
    .A2(_06823_),
    .A3(_06695_),
    .B(_06490_),
    .ZN(_06824_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13827_ (.A1(_06319_),
    .A2(_06324_),
    .A3(_06643_),
    .ZN(_06825_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13828_ (.A1(_06283_),
    .A2(_06824_),
    .B1(_06825_),
    .B2(_06642_),
    .ZN(_06826_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13829_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[29] ),
    .I1(\mod.u_arbiter.i_wb_cpu_rdt[13] ),
    .S(_06335_),
    .Z(_06827_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _13830_ (.A1(\mod.u_cpu.cpu.immdec.imm30_25[4] ),
    .A2(_06773_),
    .B1(_06812_),
    .B2(\mod.u_cpu.cpu.immdec.imm30_25[5] ),
    .C1(_06827_),
    .C2(_06339_),
    .ZN(_06828_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13831_ (.A1(_06135_),
    .A2(_06826_),
    .B(_06828_),
    .ZN(_01306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13832_ (.A1(_05790_),
    .A2(_03670_),
    .B(_03679_),
    .ZN(_06829_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13833_ (.A1(_06764_),
    .A2(_06829_),
    .ZN(_06830_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _13834_ (.A1(_06651_),
    .A2(_06829_),
    .B(_06830_),
    .C(_03682_),
    .ZN(_06831_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _13835_ (.A1(\mod.u_cpu.cpu.immdec.imm7 ),
    .A2(_03682_),
    .B(_06812_),
    .C(_06831_),
    .ZN(_06832_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13836_ (.A1(\mod.u_cpu.cpu.immdec.imm30_25[5] ),
    .A2(_06774_),
    .ZN(_06833_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13837_ (.A1(_06340_),
    .A2(_06832_),
    .A3(_06833_),
    .ZN(_01307_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _13838_ (.A1(_03331_),
    .A2(_03404_),
    .A3(_01424_),
    .B(_03334_),
    .ZN(_06834_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13839_ (.A1(_06138_),
    .A2(_06834_),
    .Z(_06835_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13840_ (.I(_06835_),
    .Z(_06836_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13841_ (.A1(_05787_),
    .A2(_06834_),
    .ZN(_06837_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13842_ (.A1(\mod.u_cpu.cpu.immdec.imm24_20[0] ),
    .A2(_06836_),
    .B1(_06837_),
    .B2(\mod.u_cpu.cpu.immdec.imm24_20[1] ),
    .ZN(_06838_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13843_ (.A1(_06677_),
    .A2(_06838_),
    .ZN(_01308_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13844_ (.A1(_06367_),
    .A2(_06743_),
    .ZN(_06839_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13845_ (.A1(_06775_),
    .A2(_06839_),
    .B(_06450_),
    .ZN(_06840_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13846_ (.A1(_06437_),
    .A2(_06662_),
    .B(_06840_),
    .ZN(_06841_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13847_ (.A1(_06803_),
    .A2(_06841_),
    .ZN(_06842_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13848_ (.A1(_06334_),
    .A2(\mod.u_arbiter.i_wb_cpu_rdt[21] ),
    .Z(_06843_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _13849_ (.A1(_06739_),
    .A2(\mod.u_arbiter.i_wb_cpu_rdt[5] ),
    .B(_06455_),
    .C(_06843_),
    .ZN(_06844_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13850_ (.A1(_06472_),
    .A2(_06443_),
    .A3(_06466_),
    .ZN(_06845_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _13851_ (.A1(_06451_),
    .A2(_06672_),
    .B(_06844_),
    .C(_06845_),
    .ZN(_06846_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13852_ (.A1(_06842_),
    .A2(_06846_),
    .B(_06483_),
    .ZN(_06847_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13853_ (.A1(\mod.u_cpu.cpu.immdec.imm24_20[1] ),
    .A2(_06836_),
    .B1(_06837_),
    .B2(\mod.u_cpu.cpu.immdec.imm24_20[2] ),
    .ZN(_06848_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13854_ (.A1(_06847_),
    .A2(_06848_),
    .ZN(_01309_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13855_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[22] ),
    .I1(\mod.u_arbiter.i_wb_cpu_rdt[6] ),
    .S(_06335_),
    .Z(_06849_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13856_ (.A1(_06397_),
    .A2(_06292_),
    .ZN(_06850_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13857_ (.A1(_06487_),
    .A2(_06850_),
    .ZN(_06851_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13858_ (.A1(_06435_),
    .A2(_06370_),
    .B(_06436_),
    .ZN(_06852_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _13859_ (.A1(_06664_),
    .A2(_06851_),
    .B1(_06852_),
    .B2(_06464_),
    .ZN(_06853_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13860_ (.A1(_06465_),
    .A2(_06744_),
    .B(_06840_),
    .ZN(_06854_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13861_ (.A1(_06853_),
    .A2(_06854_),
    .ZN(_06855_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _13862_ (.A1(_06814_),
    .A2(_06849_),
    .B(_06855_),
    .C(_06704_),
    .ZN(_06856_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13863_ (.A1(\mod.u_cpu.cpu.immdec.imm24_20[2] ),
    .A2(_06836_),
    .B1(_06837_),
    .B2(\mod.u_cpu.cpu.immdec.imm24_20[3] ),
    .ZN(_06857_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13864_ (.A1(_06856_),
    .A2(_06857_),
    .ZN(_01310_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13865_ (.A1(_06282_),
    .A2(_06294_),
    .A3(_06305_),
    .ZN(_06858_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13866_ (.A1(_06791_),
    .A2(_06672_),
    .A3(_06858_),
    .ZN(_06859_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _13867_ (.A1(_06823_),
    .A2(_06449_),
    .B(_06791_),
    .C(_06131_),
    .ZN(_06860_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13868_ (.I(_06365_),
    .Z(_06861_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _13869_ (.A1(_06694_),
    .A2(_06438_),
    .A3(_06664_),
    .A4(_06283_),
    .ZN(_06862_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13870_ (.A1(_06861_),
    .A2(_06862_),
    .ZN(_06863_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13871_ (.A1(_06840_),
    .A2(_06859_),
    .B1(_06860_),
    .B2(_06863_),
    .ZN(_06864_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _13872_ (.A1(_03503_),
    .A2(\mod.u_arbiter.i_wb_cpu_rdt[23] ),
    .Z(_06865_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13873_ (.A1(_06739_),
    .A2(\mod.u_arbiter.i_wb_cpu_rdt[7] ),
    .B(_06865_),
    .ZN(_06866_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13874_ (.A1(_06412_),
    .A2(_06834_),
    .ZN(_06867_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13875_ (.I(\mod.u_cpu.cpu.immdec.imm24_20[4] ),
    .ZN(_06868_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13876_ (.A1(_06868_),
    .A2(_06837_),
    .ZN(_06869_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13877_ (.A1(\mod.u_cpu.cpu.immdec.imm24_20[3] ),
    .A2(_06867_),
    .B(_06869_),
    .ZN(_06870_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _13878_ (.A1(_06422_),
    .A2(_06864_),
    .B1(_06866_),
    .B2(_06811_),
    .C(_06870_),
    .ZN(_01311_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13879_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[24] ),
    .I1(\mod.u_arbiter.i_wb_cpu_rdt[8] ),
    .S(_06334_),
    .Z(_06871_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13880_ (.A1(_06811_),
    .A2(_06871_),
    .ZN(_06872_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13881_ (.A1(_06426_),
    .A2(_06670_),
    .ZN(_06873_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _13882_ (.A1(_06858_),
    .A2(_06873_),
    .Z(_06874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13883_ (.A1(_06468_),
    .A2(_06874_),
    .ZN(_06875_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13884_ (.A1(_06492_),
    .A2(_06311_),
    .ZN(_06876_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _13885_ (.A1(_06735_),
    .A2(_06672_),
    .A3(_06875_),
    .A4(_06876_),
    .ZN(_06877_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13886_ (.A1(_06382_),
    .A2(_06285_),
    .B1(_06871_),
    .B2(_06441_),
    .ZN(_06878_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _13887_ (.A1(_06823_),
    .A2(_06850_),
    .B1(_06878_),
    .B2(_06423_),
    .C(_06409_),
    .ZN(_06879_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _13888_ (.A1(\mod.u_cpu.cpu.immdec.imm30_25[0] ),
    .A2(_06640_),
    .B1(_06877_),
    .B2(_06879_),
    .C(_06835_),
    .ZN(_06880_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13889_ (.A1(_06868_),
    .A2(_06836_),
    .B1(_06872_),
    .B2(_06880_),
    .ZN(_01312_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13890_ (.I(_06704_),
    .Z(_06881_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13891_ (.A1(_01426_),
    .A2(_06881_),
    .B(_06800_),
    .ZN(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13892_ (.A1(_03872_),
    .A2(_06223_),
    .ZN(_06882_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13893_ (.I0(_06578_),
    .I1(\mod.u_cpu.rf_ram.memory[112][0] ),
    .S(_06882_),
    .Z(_06883_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13894_ (.I(_06883_),
    .Z(_01314_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13895_ (.I0(_06581_),
    .I1(\mod.u_cpu.rf_ram.memory[112][1] ),
    .S(_06882_),
    .Z(_06884_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13896_ (.I(_06884_),
    .Z(_01315_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13897_ (.A1(_03342_),
    .A2(_06881_),
    .B(_06856_),
    .ZN(_01316_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13898_ (.A1(_01435_),
    .A2(_06881_),
    .B(_06847_),
    .ZN(_01317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13899_ (.A1(_01453_),
    .A2(_06140_),
    .ZN(_06885_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13900_ (.A1(_06677_),
    .A2(_06885_),
    .ZN(_01318_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13901_ (.A1(_03306_),
    .A2(_06881_),
    .B(_06689_),
    .ZN(_01319_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _13902_ (.A1(_03359_),
    .A2(_06422_),
    .B1(_06693_),
    .B2(_06463_),
    .C1(_06699_),
    .C2(_06135_),
    .ZN(_01320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13903_ (.A1(_03355_),
    .A2(_06140_),
    .ZN(_06886_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13904_ (.A1(_06707_),
    .A2(_06886_),
    .ZN(_01321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13905_ (.A1(_06481_),
    .A2(_06660_),
    .ZN(_06887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13906_ (.A1(_06065_),
    .A2(_06490_),
    .ZN(_06888_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _13907_ (.A1(_06647_),
    .A2(_06661_),
    .B1(_06682_),
    .B2(_06861_),
    .C(_06888_),
    .ZN(_06889_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13908_ (.A1(_03681_),
    .A2(_06641_),
    .B1(_06887_),
    .B2(_06889_),
    .ZN(_01322_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13909_ (.A1(_06311_),
    .A2(_06861_),
    .B1(_06443_),
    .B2(_06647_),
    .ZN(_06890_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13910_ (.A1(_03679_),
    .A2(_06649_),
    .ZN(_06891_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13911_ (.A1(_06641_),
    .A2(_06890_),
    .B(_06891_),
    .ZN(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _13912_ (.A1(_06471_),
    .A2(_06823_),
    .A3(_06390_),
    .A4(_06660_),
    .ZN(_06892_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13913_ (.A1(_06398_),
    .A2(_06452_),
    .B(_06695_),
    .ZN(_06893_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13914_ (.A1(_06476_),
    .A2(_06892_),
    .A3(_06893_),
    .ZN(_06894_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13915_ (.A1(_05790_),
    .A2(_06413_),
    .B1(_06811_),
    .B2(_06465_),
    .ZN(_06895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13916_ (.A1(_06894_),
    .A2(_06895_),
    .ZN(_01324_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13917_ (.A1(_06647_),
    .A2(_06791_),
    .B(_06640_),
    .ZN(_06896_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _13918_ (.A1(_06451_),
    .A2(_06874_),
    .B(_06487_),
    .C(_06814_),
    .ZN(_06897_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13919_ (.A1(_03403_),
    .A2(_06649_),
    .B1(_06896_),
    .B2(_06897_),
    .ZN(_06898_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _13920_ (.I(_06898_),
    .ZN(_01325_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _13921_ (.A1(_06456_),
    .A2(_06468_),
    .B1(_06861_),
    .B2(_06452_),
    .C(_06481_),
    .ZN(_06899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13922_ (.A1(_06166_),
    .A2(_06649_),
    .ZN(_06900_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13923_ (.A1(_06641_),
    .A2(_06899_),
    .B(_06900_),
    .ZN(_01326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13924_ (.A1(_04067_),
    .A2(_06030_),
    .ZN(_06901_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13925_ (.A1(_06249_),
    .A2(_06901_),
    .ZN(_06902_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13926_ (.A1(_02304_),
    .A2(_06901_),
    .B(_06902_),
    .ZN(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13927_ (.I(_06017_),
    .Z(_06903_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _13928_ (.I(_06903_),
    .Z(_06904_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _13929_ (.I0(_06904_),
    .I1(\mod.u_cpu.rf_ram.memory[111][1] ),
    .S(_06901_),
    .Z(_06905_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13930_ (.I(_06905_),
    .Z(_01328_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13931_ (.I(_05801_),
    .Z(_06906_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _13932_ (.A1(_03268_),
    .A2(\mod.u_cpu.cpu.bufreg.lsb[1] ),
    .B(_03279_),
    .C(_03269_),
    .ZN(_06907_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13933_ (.A1(_06153_),
    .A2(\mod.u_cpu.cpu.bufreg.lsb[1] ),
    .B(_03390_),
    .ZN(_06908_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _13934_ (.A1(_03394_),
    .A2(_03280_),
    .B1(_06907_),
    .B2(_06908_),
    .C(_05800_),
    .ZN(_06909_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13935_ (.I(_06909_),
    .Z(_06910_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13936_ (.I(_06910_),
    .Z(_06911_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13937_ (.I(_05792_),
    .Z(_06912_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13938_ (.A1(_05800_),
    .A2(_06909_),
    .ZN(_06913_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13939_ (.I(_06913_),
    .Z(_06914_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13940_ (.A1(_03434_),
    .A2(_06912_),
    .B(_06914_),
    .ZN(_06915_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _13941_ (.A1(_03431_),
    .A2(_06912_),
    .B(_06915_),
    .ZN(_06916_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _13942_ (.A1(_06123_),
    .A2(_06906_),
    .B1(_06911_),
    .B2(_03431_),
    .C(_06916_),
    .ZN(_01329_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13943_ (.I(_06912_),
    .Z(_06917_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13944_ (.I(_06913_),
    .Z(_06918_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13945_ (.I(_06918_),
    .Z(_06919_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13946_ (.I(_06912_),
    .Z(_06920_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13947_ (.A1(_03430_),
    .A2(_03433_),
    .Z(_06921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13948_ (.A1(_06920_),
    .A2(_06921_),
    .ZN(_06922_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _13949_ (.A1(_03438_),
    .A2(_06917_),
    .B(_06919_),
    .C(_06922_),
    .ZN(_06923_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13950_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[1] ),
    .A2(_06906_),
    .B1(_06911_),
    .B2(_03433_),
    .ZN(_06924_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13951_ (.A1(_06923_),
    .A2(_06924_),
    .ZN(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _13952_ (.A1(_03430_),
    .A2(_03433_),
    .B(_03438_),
    .ZN(_06925_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13953_ (.A1(_06920_),
    .A2(_05793_),
    .A3(_06925_),
    .ZN(_06926_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _13954_ (.A1(_03441_),
    .A2(_06917_),
    .B(_06918_),
    .C(_06926_),
    .ZN(_06927_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13955_ (.I(_06910_),
    .Z(_06928_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13956_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[2] ),
    .A2(_06906_),
    .B1(_06928_),
    .B2(_03438_),
    .ZN(_06929_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13957_ (.A1(_06927_),
    .A2(_06929_),
    .ZN(_01331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13958_ (.A1(_03441_),
    .A2(_05793_),
    .ZN(_06930_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _13959_ (.A1(_06920_),
    .A2(_05794_),
    .A3(_06930_),
    .ZN(_06931_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _13960_ (.A1(_03444_),
    .A2(_06917_),
    .B(_06918_),
    .C(_06931_),
    .ZN(_06932_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13961_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[3] ),
    .A2(_06906_),
    .B1(_06928_),
    .B2(_03441_),
    .ZN(_06933_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13962_ (.A1(_06932_),
    .A2(_06933_),
    .ZN(_01332_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _13963_ (.A1(_03444_),
    .A2(_05794_),
    .Z(_06934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13964_ (.A1(_06920_),
    .A2(_06934_),
    .ZN(_06935_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _13965_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .A2(_06917_),
    .B(_06918_),
    .C(_06935_),
    .ZN(_06936_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13966_ (.I(_05801_),
    .Z(_06937_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13967_ (.I(_06937_),
    .Z(_06938_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13968_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[4] ),
    .A2(_06938_),
    .B1(_06928_),
    .B2(_03444_),
    .ZN(_06939_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13969_ (.A1(_06936_),
    .A2(_06939_),
    .ZN(_01333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13970_ (.A1(_03412_),
    .A2(_03614_),
    .ZN(_06940_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _13971_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[5] ),
    .A2(_06940_),
    .ZN(_06941_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _13972_ (.A1(_03446_),
    .A2(_06911_),
    .B1(_06919_),
    .B2(_05798_),
    .C(_06941_),
    .ZN(_01334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13973_ (.I(_06914_),
    .Z(_06942_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13974_ (.I(_06942_),
    .Z(_06943_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13975_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[7] ),
    .A2(_06943_),
    .ZN(_06944_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13976_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[6] ),
    .A2(_06938_),
    .B1(_06928_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[6] ),
    .ZN(_06945_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13977_ (.A1(_06944_),
    .A2(_06945_),
    .ZN(_01335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13978_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[8] ),
    .A2(_06943_),
    .ZN(_06946_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13979_ (.I(_06910_),
    .Z(_06947_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13980_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[7] ),
    .A2(_06938_),
    .B1(_06947_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[7] ),
    .ZN(_06948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13981_ (.A1(_06946_),
    .A2(_06948_),
    .ZN(_01336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13982_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[9] ),
    .A2(_06943_),
    .ZN(_06949_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13983_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[8] ),
    .A2(_06938_),
    .B1(_06947_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[8] ),
    .ZN(_06950_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13984_ (.A1(_06949_),
    .A2(_06950_),
    .ZN(_01337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13985_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[10] ),
    .A2(_06943_),
    .ZN(_06951_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13986_ (.I(_06937_),
    .Z(_06952_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13987_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[9] ),
    .A2(_06952_),
    .B1(_06947_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[9] ),
    .ZN(_06953_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13988_ (.A1(_06951_),
    .A2(_06953_),
    .ZN(_01338_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13989_ (.I(_06942_),
    .Z(_06954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13990_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[11] ),
    .A2(_06954_),
    .ZN(_06955_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13991_ (.A1(_03449_),
    .A2(_06952_),
    .B1(_06947_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[10] ),
    .ZN(_06956_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13992_ (.A1(_06955_),
    .A2(_06956_),
    .ZN(_01339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13993_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[12] ),
    .A2(_06954_),
    .ZN(_06957_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _13994_ (.I(_06910_),
    .Z(_06958_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13995_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[11] ),
    .A2(_06952_),
    .B1(_06958_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[11] ),
    .ZN(_06959_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13996_ (.A1(_06957_),
    .A2(_06959_),
    .ZN(_01340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13997_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[13] ),
    .A2(_06954_),
    .ZN(_06960_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _13998_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[12] ),
    .A2(_06952_),
    .B1(_06958_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[12] ),
    .ZN(_06961_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _13999_ (.A1(_06960_),
    .A2(_06961_),
    .ZN(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14000_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[14] ),
    .A2(_06954_),
    .ZN(_06962_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14001_ (.I(_05801_),
    .Z(_06963_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14002_ (.I(_06963_),
    .Z(_06964_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _14003_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[13] ),
    .A2(_06964_),
    .B1(_06958_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[13] ),
    .ZN(_06965_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14004_ (.A1(_06962_),
    .A2(_06965_),
    .ZN(_01342_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14005_ (.I(_06942_),
    .Z(_06966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14006_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[15] ),
    .A2(_06966_),
    .ZN(_06967_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _14007_ (.A1(_03456_),
    .A2(_06964_),
    .B1(_06958_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[14] ),
    .ZN(_06968_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14008_ (.A1(_06967_),
    .A2(_06968_),
    .ZN(_01343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14009_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[16] ),
    .A2(_06966_),
    .ZN(_06969_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14010_ (.I(_06909_),
    .Z(_06970_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14011_ (.I(_06970_),
    .Z(_06971_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _14012_ (.A1(_03458_),
    .A2(_06964_),
    .B1(_06971_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[15] ),
    .ZN(_06972_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14013_ (.A1(_06969_),
    .A2(_06972_),
    .ZN(_01344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14014_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[17] ),
    .A2(_06966_),
    .ZN(_06973_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _14015_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[16] ),
    .A2(_06964_),
    .B1(_06971_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[16] ),
    .ZN(_06974_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14016_ (.A1(_06973_),
    .A2(_06974_),
    .ZN(_01345_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14017_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[18] ),
    .A2(_06966_),
    .ZN(_06975_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14018_ (.I(_06963_),
    .Z(_06976_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _14019_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[17] ),
    .A2(_06976_),
    .B1(_06971_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[17] ),
    .ZN(_06977_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14020_ (.A1(_06975_),
    .A2(_06977_),
    .ZN(_01346_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14021_ (.I(_06942_),
    .Z(_06978_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14022_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[19] ),
    .A2(_06978_),
    .ZN(_06979_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _14023_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[18] ),
    .A2(_06976_),
    .B1(_06971_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[18] ),
    .ZN(_06980_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14024_ (.A1(_06979_),
    .A2(_06980_),
    .ZN(_01347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14025_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[20] ),
    .A2(_06978_),
    .ZN(_06981_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14026_ (.I(_06970_),
    .Z(_06982_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _14027_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[19] ),
    .A2(_06976_),
    .B1(_06982_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[19] ),
    .ZN(_06983_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14028_ (.A1(_06981_),
    .A2(_06983_),
    .ZN(_01348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14029_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[21] ),
    .A2(_06978_),
    .ZN(_06984_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _14030_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[20] ),
    .A2(_06976_),
    .B1(_06982_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[20] ),
    .ZN(_06985_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14031_ (.A1(_06984_),
    .A2(_06985_),
    .ZN(_01349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14032_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[22] ),
    .A2(_06978_),
    .ZN(_06986_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14033_ (.I(_06963_),
    .Z(_06987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _14034_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[21] ),
    .A2(_06987_),
    .B1(_06982_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[21] ),
    .ZN(_06988_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14035_ (.A1(_06986_),
    .A2(_06988_),
    .ZN(_01350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14036_ (.I(_06914_),
    .Z(_06989_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14037_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[23] ),
    .A2(_06989_),
    .ZN(_06990_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _14038_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[22] ),
    .A2(_06987_),
    .B1(_06982_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[22] ),
    .ZN(_06991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14039_ (.A1(_06990_),
    .A2(_06991_),
    .ZN(_01351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14040_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[24] ),
    .A2(_06989_),
    .ZN(_06992_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14041_ (.I(_06970_),
    .Z(_06993_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _14042_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[23] ),
    .A2(_06987_),
    .B1(_06993_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[23] ),
    .ZN(_06994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14043_ (.A1(_06992_),
    .A2(_06994_),
    .ZN(_01352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14044_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[25] ),
    .A2(_06989_),
    .ZN(_06995_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _14045_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[24] ),
    .A2(_06987_),
    .B1(_06993_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[24] ),
    .ZN(_06996_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14046_ (.A1(_06995_),
    .A2(_06996_),
    .ZN(_01353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14047_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[26] ),
    .A2(_06989_),
    .ZN(_06997_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14048_ (.I(_06963_),
    .Z(_06998_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _14049_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[25] ),
    .A2(_06998_),
    .B1(_06993_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[25] ),
    .ZN(_06999_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14050_ (.A1(_06997_),
    .A2(_06999_),
    .ZN(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14051_ (.I(_06914_),
    .Z(_07000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14052_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[27] ),
    .A2(_07000_),
    .ZN(_07001_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _14053_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[26] ),
    .A2(_06998_),
    .B1(_06993_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[26] ),
    .ZN(_07002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14054_ (.A1(_07001_),
    .A2(_07002_),
    .ZN(_01355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14055_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[28] ),
    .A2(_07000_),
    .ZN(_07003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14056_ (.I(_06970_),
    .Z(_07004_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _14057_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[27] ),
    .A2(_06998_),
    .B1(_07004_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[27] ),
    .ZN(_07005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14058_ (.A1(_07003_),
    .A2(_07005_),
    .ZN(_01356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14059_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[29] ),
    .A2(_07000_),
    .ZN(_07006_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _14060_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[28] ),
    .A2(_06998_),
    .B1(_07004_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[28] ),
    .ZN(_07007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14061_ (.A1(_07006_),
    .A2(_07007_),
    .ZN(_01357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14062_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[30] ),
    .A2(_07000_),
    .ZN(_07008_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _14063_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[29] ),
    .A2(_06937_),
    .B1(_07004_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[29] ),
    .ZN(_07009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14064_ (.A1(_07008_),
    .A2(_07009_),
    .ZN(_01358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14065_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[31] ),
    .A2(_06919_),
    .ZN(_07010_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _14066_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[30] ),
    .A2(_06937_),
    .B1(_07004_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[30] ),
    .ZN(_07011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14067_ (.A1(_07010_),
    .A2(_07011_),
    .ZN(_01359_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14068_ (.I(_03309_),
    .ZN(_07012_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14069_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[31] ),
    .A2(_06940_),
    .ZN(_07013_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _14070_ (.A1(_03483_),
    .A2(_06911_),
    .B1(_06919_),
    .B2(_07012_),
    .C(_07013_),
    .ZN(_01360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14071_ (.I(_05630_),
    .Z(_07014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14072_ (.A1(_03858_),
    .A2(_07014_),
    .ZN(_07015_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14073_ (.I0(_06578_),
    .I1(\mod.u_cpu.rf_ram.memory[114][0] ),
    .S(_07015_),
    .Z(_07016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14074_ (.I(_07016_),
    .Z(_01361_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14075_ (.I0(_06904_),
    .I1(\mod.u_cpu.rf_ram.memory[114][1] ),
    .S(_07015_),
    .Z(_07017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14076_ (.I(_07017_),
    .Z(_01362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14077_ (.A1(_03910_),
    .A2(_04996_),
    .ZN(_07018_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14078_ (.I0(_06578_),
    .I1(\mod.u_cpu.rf_ram.memory[299][0] ),
    .S(_07018_),
    .Z(_07019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14079_ (.I(_07019_),
    .Z(_01363_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14080_ (.I0(_06904_),
    .I1(\mod.u_cpu.rf_ram.memory[299][1] ),
    .S(_07018_),
    .Z(_07020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14081_ (.I(_07020_),
    .Z(_01364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14082_ (.I(_06577_),
    .Z(_07021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14083_ (.A1(_03865_),
    .A2(_07014_),
    .ZN(_07022_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14084_ (.I0(_07021_),
    .I1(\mod.u_cpu.rf_ram.memory[113][0] ),
    .S(_07022_),
    .Z(_07023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14085_ (.I(_07023_),
    .Z(_01365_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14086_ (.I0(_06904_),
    .I1(\mod.u_cpu.rf_ram.memory[113][1] ),
    .S(_07022_),
    .Z(_07024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14087_ (.I(_07024_),
    .Z(_01366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14088_ (.A1(_03836_),
    .A2(_05279_),
    .ZN(_07025_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14089_ (.I(_03774_),
    .Z(_07026_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14090_ (.A1(_07026_),
    .A2(_07025_),
    .ZN(_07027_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14091_ (.A1(_02258_),
    .A2(_07025_),
    .B(_07027_),
    .ZN(_01367_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14092_ (.I(_06903_),
    .Z(_07028_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14093_ (.I0(_07028_),
    .I1(\mod.u_cpu.rf_ram.memory[245][1] ),
    .S(_07025_),
    .Z(_07029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14094_ (.I(_07029_),
    .Z(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14095_ (.A1(_03804_),
    .A2(_07014_),
    .ZN(_07030_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14096_ (.I0(_07021_),
    .I1(\mod.u_cpu.rf_ram.memory[120][0] ),
    .S(_07030_),
    .Z(_07031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14097_ (.I(_07031_),
    .Z(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14098_ (.I0(_07028_),
    .I1(\mod.u_cpu.rf_ram.memory[120][1] ),
    .S(_07030_),
    .Z(_07032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14099_ (.I(_07032_),
    .Z(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14100_ (.A1(_03885_),
    .A2(_07014_),
    .ZN(_07033_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14101_ (.I0(_07021_),
    .I1(\mod.u_cpu.rf_ram.memory[110][0] ),
    .S(_07033_),
    .Z(_07034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14102_ (.I(_07034_),
    .Z(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14103_ (.I0(_07028_),
    .I1(\mod.u_cpu.rf_ram.memory[110][1] ),
    .S(_07033_),
    .Z(_07035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14104_ (.I(_07035_),
    .Z(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14105_ (.A1(_03836_),
    .A2(_05720_),
    .ZN(_07036_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14106_ (.A1(_07026_),
    .A2(_07036_),
    .ZN(_07037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14107_ (.A1(_02326_),
    .A2(_07036_),
    .B(_07037_),
    .ZN(_01373_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14108_ (.I0(_07028_),
    .I1(\mod.u_cpu.rf_ram.memory[117][1] ),
    .S(_07036_),
    .Z(_07038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14109_ (.I(_07038_),
    .Z(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14110_ (.A1(_03823_),
    .A2(_05397_),
    .ZN(_07039_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14111_ (.I0(_07021_),
    .I1(\mod.u_cpu.rf_ram.memory[87][0] ),
    .S(_07039_),
    .Z(_07040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14112_ (.I(_07040_),
    .Z(_01375_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14113_ (.I(_06903_),
    .Z(_07041_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14114_ (.I0(_07041_),
    .I1(\mod.u_cpu.rf_ram.memory[87][1] ),
    .S(_07039_),
    .Z(_07042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14115_ (.I(_07042_),
    .Z(_01376_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14116_ (.I(_06577_),
    .Z(_07043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14117_ (.A1(_06181_),
    .A2(_03911_),
    .ZN(_07044_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14118_ (.I0(_07043_),
    .I1(\mod.u_cpu.rf_ram.memory[11][0] ),
    .S(_07044_),
    .Z(_07045_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14119_ (.I(_07045_),
    .Z(_01377_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14120_ (.I0(_07041_),
    .I1(\mod.u_cpu.rf_ram.memory[11][1] ),
    .S(_07044_),
    .Z(_07046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14121_ (.I(_07046_),
    .Z(_01378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14122_ (.A1(_03842_),
    .A2(_05631_),
    .ZN(_07047_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14123_ (.I0(_07043_),
    .I1(\mod.u_cpu.rf_ram.memory[116][0] ),
    .S(_07047_),
    .Z(_07048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14124_ (.I(_07048_),
    .Z(_01379_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14125_ (.I0(_07041_),
    .I1(\mod.u_cpu.rf_ram.memory[116][1] ),
    .S(_07047_),
    .Z(_07049_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14126_ (.I(_07049_),
    .Z(_01380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14127_ (.A1(_03828_),
    .A2(_05631_),
    .ZN(_07050_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14128_ (.I0(_07043_),
    .I1(\mod.u_cpu.rf_ram.memory[118][0] ),
    .S(_07050_),
    .Z(_07051_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14129_ (.I(_07051_),
    .Z(_01381_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14130_ (.I0(_07041_),
    .I1(\mod.u_cpu.rf_ram.memory[118][1] ),
    .S(_07050_),
    .Z(_07052_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14131_ (.I(_07052_),
    .Z(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14132_ (.A1(_03850_),
    .A2(_05631_),
    .ZN(_07053_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14133_ (.I0(_07043_),
    .I1(\mod.u_cpu.rf_ram.memory[115][0] ),
    .S(_07053_),
    .Z(_07054_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14134_ (.I(_07054_),
    .Z(_01383_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14135_ (.I(_06903_),
    .Z(_07055_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14136_ (.I0(_07055_),
    .I1(\mod.u_cpu.rf_ram.memory[115][1] ),
    .S(_07053_),
    .Z(_07056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14137_ (.I(_07056_),
    .Z(_01384_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14138_ (.I(_06577_),
    .Z(_07057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14139_ (.A1(_03980_),
    .A2(_04996_),
    .ZN(_07058_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14140_ (.I0(_07057_),
    .I1(\mod.u_cpu.rf_ram.memory[289][0] ),
    .S(_07058_),
    .Z(_07059_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14141_ (.I(_07059_),
    .Z(_01385_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14142_ (.I0(_07055_),
    .I1(\mod.u_cpu.rf_ram.memory[289][1] ),
    .S(_07058_),
    .Z(_07060_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14143_ (.I(_07060_),
    .Z(_01386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14144_ (.A1(_03796_),
    .A2(_05397_),
    .ZN(_07061_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14145_ (.I0(_07057_),
    .I1(\mod.u_cpu.rf_ram.memory[90][0] ),
    .S(_07061_),
    .Z(_07062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14146_ (.I(_07062_),
    .Z(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14147_ (.I0(_07055_),
    .I1(\mod.u_cpu.rf_ram.memory[90][1] ),
    .S(_07061_),
    .Z(_07063_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14148_ (.I(_07063_),
    .Z(_01388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14149_ (.A1(_03822_),
    .A2(_05254_),
    .ZN(_07064_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14150_ (.A1(_07026_),
    .A2(_07064_),
    .ZN(_07065_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14151_ (.A1(_02261_),
    .A2(_07064_),
    .B(_07065_),
    .ZN(_01389_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14152_ (.I0(_07055_),
    .I1(\mod.u_cpu.rf_ram.memory[247][1] ),
    .S(_07064_),
    .Z(_07066_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14153_ (.I(_07066_),
    .Z(_01390_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14154_ (.I(_06063_),
    .ZN(_07067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14155_ (.A1(_06057_),
    .A2(_06111_),
    .ZN(_07068_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14156_ (.A1(_07067_),
    .A2(_03284_),
    .B(_07068_),
    .ZN(_01391_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14157_ (.A1(_06056_),
    .A2(\mod.u_cpu.cpu.state.o_cnt_r[2] ),
    .Z(_07069_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14158_ (.I(_07069_),
    .Z(_01407_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _14159_ (.A1(_06153_),
    .A2(_03270_),
    .A3(_01407_),
    .Z(_07070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14160_ (.I(_07070_),
    .Z(_01392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14161_ (.A1(_07067_),
    .A2(\mod.u_cpu.cpu.ctrl.i_jump ),
    .ZN(_07071_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14162_ (.A1(_03363_),
    .A2(_06631_),
    .Z(_07072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14163_ (.A1(_06062_),
    .A2(_06568_),
    .ZN(_07073_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14164_ (.A1(_03298_),
    .A2(_07073_),
    .ZN(_07074_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14165_ (.A1(_03670_),
    .A2(_07072_),
    .B(_07074_),
    .ZN(_07075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14166_ (.I(_06046_),
    .Z(_07076_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14167_ (.A1(_07071_),
    .A2(_07075_),
    .B(_07076_),
    .ZN(_01393_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _14168_ (.A1(_05790_),
    .A2(_06166_),
    .A3(_03393_),
    .A4(_07073_),
    .ZN(_07077_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14169_ (.A1(_05780_),
    .A2(_07067_),
    .B(_07077_),
    .ZN(_07078_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14170_ (.A1(_06047_),
    .A2(_07078_),
    .ZN(_01395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14171_ (.A1(_03804_),
    .A2(_05397_),
    .ZN(_07079_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14172_ (.I0(_07057_),
    .I1(\mod.u_cpu.rf_ram.memory[88][0] ),
    .S(_07079_),
    .Z(_07080_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14173_ (.I(_07080_),
    .Z(_01396_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _14174_ (.I(_03928_),
    .Z(_07081_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14175_ (.I0(_07081_),
    .I1(\mod.u_cpu.rf_ram.memory[88][1] ),
    .S(_07079_),
    .Z(_07082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14176_ (.I(_07082_),
    .Z(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14177_ (.A1(_06181_),
    .A2(_03933_),
    .ZN(_07083_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14178_ (.I0(_07057_),
    .I1(\mod.u_cpu.rf_ram.memory[8][0] ),
    .S(_07083_),
    .Z(_07084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14179_ (.I(_07084_),
    .Z(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14180_ (.I0(_07081_),
    .I1(\mod.u_cpu.rf_ram.memory[8][1] ),
    .S(_07083_),
    .Z(_07085_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14181_ (.I(_07085_),
    .Z(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14182_ (.A1(_03822_),
    .A2(_05124_),
    .ZN(_07086_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14183_ (.A1(_07026_),
    .A2(_07086_),
    .ZN(_07087_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14184_ (.A1(_01985_),
    .A2(_07086_),
    .B(_07087_),
    .ZN(_01400_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14185_ (.I0(_07081_),
    .I1(\mod.u_cpu.rf_ram.memory[279][1] ),
    .S(_07086_),
    .Z(_07088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14186_ (.I(_07088_),
    .Z(_01401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14187_ (.A1(_03842_),
    .A2(_05263_),
    .ZN(_07089_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14188_ (.I0(_03699_),
    .I1(\mod.u_cpu.rf_ram.memory[244][0] ),
    .S(_07089_),
    .Z(_07090_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14189_ (.I(_07090_),
    .Z(_01402_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14190_ (.I0(_07081_),
    .I1(\mod.u_cpu.rf_ram.memory[244][1] ),
    .S(_07089_),
    .Z(_07091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14191_ (.I(_07091_),
    .Z(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _14192_ (.I(\mod.u_cpu.rf_ram_if.rgnt ),
    .ZN(_07092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14193_ (.A1(_07092_),
    .A2(_05803_),
    .ZN(_07093_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _14194_ (.A1(_07067_),
    .A2(_03389_),
    .B1(_03674_),
    .B2(_07093_),
    .ZN(_07094_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14195_ (.A1(_07076_),
    .A2(_07094_),
    .ZN(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _14196_ (.A1(_06057_),
    .A2(_03388_),
    .Z(_07095_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14197_ (.I(_07095_),
    .Z(_01405_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14198_ (.A1(_07076_),
    .A2(_03320_),
    .ZN(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14199_ (.A1(_03389_),
    .A2(\mod.u_cpu.cpu.state.o_cnt[2] ),
    .ZN(_07096_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _14200_ (.A1(_06046_),
    .A2(_06151_),
    .A3(_07096_),
    .ZN(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14201_ (.A1(_06152_),
    .A2(_06151_),
    .B(_06056_),
    .ZN(_07097_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _14202_ (.A1(_06152_),
    .A2(_06151_),
    .B(_07097_),
    .ZN(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14203_ (.A1(_06152_),
    .A2(_06150_),
    .ZN(_07098_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _14204_ (.A1(_06153_),
    .A2(_07098_),
    .Z(_07099_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14205_ (.A1(_07076_),
    .A2(_07099_),
    .ZN(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _14206_ (.A1(_06047_),
    .A2(_07073_),
    .ZN(_01411_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _14207_ (.A1(_03895_),
    .A2(_05210_),
    .ZN(_07100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14208_ (.A1(_03775_),
    .A2(_07100_),
    .ZN(_07101_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _14209_ (.A1(_02023_),
    .A2(_07100_),
    .B(_07101_),
    .ZN(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14210_ (.I0(\mod.u_cpu.rf_ram.memory[269][1] ),
    .I1(_06221_),
    .S(_07100_),
    .Z(_07102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14211_ (.I(_07102_),
    .Z(_01413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14212_ (.A1(_03968_),
    .A2(_05120_),
    .ZN(_07103_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14213_ (.I0(_03699_),
    .I1(\mod.u_cpu.rf_ram.memory[259][0] ),
    .S(_07103_),
    .Z(_07104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14214_ (.I(_07104_),
    .Z(_01414_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14215_ (.I0(_03735_),
    .I1(\mod.u_cpu.rf_ram.memory[259][1] ),
    .S(_07103_),
    .Z(_07105_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14216_ (.I(_07105_),
    .Z(_01415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _14217_ (.A1(_04025_),
    .A2(_05263_),
    .ZN(_07106_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14218_ (.I0(_03699_),
    .I1(\mod.u_cpu.rf_ram.memory[249][0] ),
    .S(_07106_),
    .Z(_07107_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14219_ (.I(_07107_),
    .Z(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _14220_ (.I0(_03735_),
    .I1(\mod.u_cpu.rf_ram.memory[249][1] ),
    .S(_07106_),
    .Z(_07108_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _14221_ (.I(_07108_),
    .Z(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14222_ (.D(_00078_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14223_ (.D(_00079_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14224_ (.D(_00000_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.rdata[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14225_ (.D(_00001_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.rdata[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14226_ (.D(_00080_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[574][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14227_ (.D(_00081_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[574][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14228_ (.D(_00082_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[573][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14229_ (.D(_00083_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[573][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14230_ (.D(_00084_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[572][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14231_ (.D(_00085_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[572][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14232_ (.D(_00086_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[571][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14233_ (.D(_00087_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[571][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14234_ (.D(_00088_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[570][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14235_ (.D(_00089_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[570][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14236_ (.D(_00090_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[56][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14237_ (.D(_00091_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[56][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14238_ (.D(_00092_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[568][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14239_ (.D(_00093_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[568][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14240_ (.D(_00094_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[567][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14241_ (.D(_00095_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[567][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14242_ (.D(_00096_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[566][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14243_ (.D(_00097_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[566][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14244_ (.D(_00098_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[565][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14245_ (.D(_00099_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[565][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14246_ (.D(_00100_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[564][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14247_ (.D(_00101_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[564][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14248_ (.D(_00102_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[563][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14249_ (.D(_00103_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[563][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14250_ (.D(_00104_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[562][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14251_ (.D(_00105_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[562][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14252_ (.D(_00106_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[561][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14253_ (.D(_00107_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[561][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14254_ (.D(_00108_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[560][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14255_ (.D(_00109_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[560][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14256_ (.D(_00110_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[55][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14257_ (.D(_00111_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[55][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14258_ (.D(_00112_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[558][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14259_ (.D(_00113_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[558][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14260_ (.D(_00114_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[557][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14261_ (.D(_00115_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[557][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14262_ (.D(_00116_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[556][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14263_ (.D(_00117_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[556][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14264_ (.D(_00118_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[555][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14265_ (.D(_00119_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[555][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14266_ (.D(_00120_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[554][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14267_ (.D(_00121_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[554][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14268_ (.D(_00122_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[553][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14269_ (.D(_00123_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[553][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14270_ (.D(_00124_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[552][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14271_ (.D(_00125_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[552][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14272_ (.D(_00126_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[551][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14273_ (.D(_00127_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[551][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14274_ (.D(_00128_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[550][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14275_ (.D(_00129_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[550][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14276_ (.D(_00130_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[54][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14277_ (.D(_00131_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[54][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14278_ (.D(_00132_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[548][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14279_ (.D(_00133_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[548][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14280_ (.D(_00134_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[547][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14281_ (.D(_00135_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[547][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14282_ (.D(_00136_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[546][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14283_ (.D(_00137_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[546][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14284_ (.D(_00138_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[545][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14285_ (.D(_00139_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[545][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14286_ (.D(_00140_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[544][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14287_ (.D(_00141_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[544][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14288_ (.D(_00142_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[543][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14289_ (.D(_00143_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[543][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14290_ (.D(_00144_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[542][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14291_ (.D(_00145_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[542][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14292_ (.D(_00146_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[541][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14293_ (.D(_00147_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[541][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14294_ (.D(_00148_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[540][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14295_ (.D(_00149_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[540][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14296_ (.D(_00150_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[53][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14297_ (.D(_00151_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[53][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14298_ (.D(_00152_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[538][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14299_ (.D(_00153_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[538][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14300_ (.D(_00154_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[537][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14301_ (.D(_00155_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[537][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14302_ (.D(_00156_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[536][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14303_ (.D(_00157_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[536][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14304_ (.D(_00158_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[535][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14305_ (.D(_00159_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[535][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14306_ (.D(_00160_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[534][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14307_ (.D(_00161_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[534][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14308_ (.D(_00162_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[533][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14309_ (.D(_00163_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[533][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14310_ (.D(_00164_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[532][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14311_ (.D(_00165_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[532][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14312_ (.D(_00166_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[531][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14313_ (.D(_00167_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[531][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14314_ (.D(_00168_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[530][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14315_ (.D(_00169_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[530][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14316_ (.D(_00170_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[52][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14317_ (.D(_00171_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[52][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14318_ (.D(_00172_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[528][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14319_ (.D(_00173_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[528][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14320_ (.D(_00174_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[527][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14321_ (.D(_00175_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[527][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14322_ (.D(_00176_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[526][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14323_ (.D(_00177_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[526][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14324_ (.D(_00178_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[525][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14325_ (.D(_00179_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[525][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14326_ (.D(_00180_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[524][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14327_ (.D(_00181_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[524][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14328_ (.D(_00182_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[523][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14329_ (.D(_00183_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[523][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14330_ (.D(_00184_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[522][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14331_ (.D(_00185_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[522][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14332_ (.D(_00186_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[521][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14333_ (.D(_00187_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[521][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14334_ (.D(_00188_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[520][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14335_ (.D(_00189_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[520][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14336_ (.D(_00190_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[51][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14337_ (.D(_00191_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[51][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14338_ (.D(_00192_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[518][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14339_ (.D(_00193_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[518][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14340_ (.D(_00194_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[517][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14341_ (.D(_00195_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[517][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14342_ (.D(_00196_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[516][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14343_ (.D(_00197_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[516][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14344_ (.D(_00198_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[515][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14345_ (.D(_00199_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[515][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14346_ (.D(_00200_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[514][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14347_ (.D(_00201_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[514][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14348_ (.D(_00202_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[513][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14349_ (.D(_00203_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[513][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14350_ (.D(_00204_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[512][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14351_ (.D(_00205_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[512][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14352_ (.D(_00206_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[511][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14353_ (.D(_00207_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[511][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14354_ (.D(_00208_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[510][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14355_ (.D(_00209_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[510][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14356_ (.D(_00210_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[50][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14357_ (.D(_00211_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[50][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14358_ (.D(_00212_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[508][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14359_ (.D(_00213_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[508][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14360_ (.D(_00214_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[507][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14361_ (.D(_00215_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[507][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14362_ (.D(_00216_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[506][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14363_ (.D(_00217_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[506][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14364_ (.D(_00218_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[505][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14365_ (.D(_00219_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[505][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14366_ (.D(_00220_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[504][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14367_ (.D(_00221_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[504][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14368_ (.D(_00222_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[503][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14369_ (.D(_00223_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[503][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14370_ (.D(_00224_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[502][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14371_ (.D(_00225_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[502][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14372_ (.D(_00226_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[501][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14373_ (.D(_00227_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[501][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14374_ (.D(_00228_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[500][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14375_ (.D(_00229_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[500][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14376_ (.D(_00230_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14377_ (.D(_00231_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14378_ (.D(_00232_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[498][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14379_ (.D(_00233_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[498][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14380_ (.D(_00234_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[497][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14381_ (.D(_00235_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[497][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14382_ (.D(_00236_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[496][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14383_ (.D(_00237_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[496][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14384_ (.D(_00238_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[495][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14385_ (.D(_00239_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[495][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14386_ (.D(_00240_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[494][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14387_ (.D(_00241_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[494][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14388_ (.D(_00242_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[493][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14389_ (.D(_00243_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[493][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14390_ (.D(_00244_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[492][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14391_ (.D(_00245_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[492][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14392_ (.D(_00246_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[491][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14393_ (.D(_00247_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[491][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14394_ (.D(_00248_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[490][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14395_ (.D(_00249_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[490][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14396_ (.D(_00250_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[48][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14397_ (.D(_00251_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[48][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14398_ (.D(_00252_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[488][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14399_ (.D(_00253_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[488][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14400_ (.D(_00254_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[487][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14401_ (.D(_00255_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[487][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14402_ (.D(_00256_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[486][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14403_ (.D(_00257_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[486][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14404_ (.D(_00258_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[485][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14405_ (.D(_00259_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[485][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14406_ (.D(_00260_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[484][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14407_ (.D(_00261_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[484][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14408_ (.D(_00262_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[483][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14409_ (.D(_00263_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[483][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14410_ (.D(_00264_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[482][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14411_ (.D(_00265_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[482][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14412_ (.D(_00266_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[481][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14413_ (.D(_00267_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[481][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14414_ (.D(_00268_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[480][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14415_ (.D(_00269_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[480][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14416_ (.D(_00270_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[47][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14417_ (.D(_00271_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[47][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14418_ (.D(_00272_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[478][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14419_ (.D(_00273_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[478][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14420_ (.D(_00274_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[477][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14421_ (.D(_00275_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[477][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14422_ (.D(_00276_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[476][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14423_ (.D(_00277_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[476][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14424_ (.D(_00278_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[475][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14425_ (.D(_00279_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[475][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14426_ (.D(_00280_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[474][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14427_ (.D(_00281_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[474][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14428_ (.D(_00282_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[473][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14429_ (.D(_00283_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[473][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14430_ (.D(_00284_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[472][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14431_ (.D(_00285_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[472][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14432_ (.D(_00286_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[471][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14433_ (.D(_00287_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[471][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14434_ (.D(_00288_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[470][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14435_ (.D(_00289_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[470][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14436_ (.D(_00290_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[46][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14437_ (.D(_00291_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[46][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14438_ (.D(_00292_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[468][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14439_ (.D(_00293_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[468][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14440_ (.D(_00294_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[467][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14441_ (.D(_00295_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[467][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14442_ (.D(_00296_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[466][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14443_ (.D(_00297_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[466][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14444_ (.D(_00298_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[465][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14445_ (.D(_00299_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[465][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14446_ (.D(_00300_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[464][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14447_ (.D(_00301_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[464][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14448_ (.D(_00302_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[463][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14449_ (.D(_00303_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[463][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14450_ (.D(_00304_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[462][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14451_ (.D(_00305_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[462][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14452_ (.D(_00306_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[461][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14453_ (.D(_00307_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[461][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14454_ (.D(_00308_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[460][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14455_ (.D(_00309_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[460][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14456_ (.D(_00310_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[45][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14457_ (.D(_00311_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[45][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14458_ (.D(_00312_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[458][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14459_ (.D(_00313_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[458][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14460_ (.D(_00314_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[457][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14461_ (.D(_00315_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[457][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14462_ (.D(_00316_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[456][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14463_ (.D(_00317_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[456][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14464_ (.D(_00318_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[455][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14465_ (.D(_00319_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[455][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14466_ (.D(_00320_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[454][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14467_ (.D(_00321_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[454][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14468_ (.D(_00322_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[453][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14469_ (.D(_00323_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[453][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14470_ (.D(_00324_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[452][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14471_ (.D(_00325_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[452][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14472_ (.D(_00326_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[451][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14473_ (.D(_00327_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[451][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14474_ (.D(_00328_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[450][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14475_ (.D(_00329_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[450][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14476_ (.D(_00330_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[44][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14477_ (.D(_00331_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[44][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14478_ (.D(_00332_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[448][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14479_ (.D(_00333_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[448][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14480_ (.D(_00334_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[447][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14481_ (.D(_00335_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[447][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14482_ (.D(_00336_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[446][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14483_ (.D(_00337_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[446][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14484_ (.D(_00338_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[445][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14485_ (.D(_00339_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[445][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14486_ (.D(_00340_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[444][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14487_ (.D(_00341_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[444][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14488_ (.D(_00342_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[443][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14489_ (.D(_00343_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[443][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14490_ (.D(_00344_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[442][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14491_ (.D(_00345_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[442][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14492_ (.D(_00346_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[441][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14493_ (.D(_00347_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[441][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14494_ (.D(_00348_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[440][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14495_ (.D(_00349_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[440][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14496_ (.D(_00350_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[43][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14497_ (.D(_00351_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[43][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14498_ (.D(_00352_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[438][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14499_ (.D(_00353_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[438][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14500_ (.D(_00354_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[437][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14501_ (.D(_00355_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[437][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14502_ (.D(_00356_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[436][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14503_ (.D(_00357_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[436][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14504_ (.D(_00358_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[435][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14505_ (.D(_00359_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[435][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14506_ (.D(_00360_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[434][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14507_ (.D(_00361_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[434][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14508_ (.D(_00362_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[433][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14509_ (.D(_00363_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[433][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14510_ (.D(_00364_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[432][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14511_ (.D(_00365_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[432][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14512_ (.D(_00366_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[431][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14513_ (.D(_00367_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[431][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14514_ (.D(_00368_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[430][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14515_ (.D(_00369_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[430][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14516_ (.D(_00370_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[42][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14517_ (.D(_00371_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[42][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14518_ (.D(_00372_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[428][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14519_ (.D(_00373_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[428][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14520_ (.D(_00374_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[427][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14521_ (.D(_00375_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[427][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14522_ (.D(_00376_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[426][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14523_ (.D(_00377_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[426][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14524_ (.D(_00378_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[425][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14525_ (.D(_00379_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[425][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14526_ (.D(_00380_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[424][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14527_ (.D(_00381_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[424][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14528_ (.D(_00382_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[423][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14529_ (.D(_00383_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[423][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14530_ (.D(_00384_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[422][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14531_ (.D(_00385_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[422][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14532_ (.D(_00386_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[421][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14533_ (.D(_00387_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[421][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14534_ (.D(_00388_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[420][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14535_ (.D(_00389_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[420][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14536_ (.D(_00390_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[41][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14537_ (.D(_00391_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[41][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14538_ (.D(_00392_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[418][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14539_ (.D(_00393_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[418][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14540_ (.D(_00394_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[417][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14541_ (.D(_00395_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[417][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14542_ (.D(_00396_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[416][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14543_ (.D(_00397_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[416][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14544_ (.D(_00398_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[415][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14545_ (.D(_00399_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[415][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14546_ (.D(_00400_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[414][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14547_ (.D(_00401_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[414][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14548_ (.D(_00402_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[413][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14549_ (.D(_00403_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[413][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14550_ (.D(_00404_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[412][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14551_ (.D(_00405_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[412][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14552_ (.D(_00406_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[411][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14553_ (.D(_00407_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[411][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14554_ (.D(_00408_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[410][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14555_ (.D(_00409_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[410][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14556_ (.D(_00410_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[40][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14557_ (.D(_00411_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[40][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14558_ (.D(_00412_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[408][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14559_ (.D(_00413_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[408][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14560_ (.D(_00414_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[407][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14561_ (.D(_00415_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[407][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14562_ (.D(_00416_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[406][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14563_ (.D(_00417_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[406][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14564_ (.D(_00418_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[405][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14565_ (.D(_00419_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[405][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14566_ (.D(_00420_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[404][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14567_ (.D(_00421_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[404][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14568_ (.D(_00422_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[403][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14569_ (.D(_00423_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[403][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14570_ (.D(_00424_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[402][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14571_ (.D(_00425_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[402][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14572_ (.D(_00426_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[401][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14573_ (.D(_00427_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[401][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14574_ (.D(_00428_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[400][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14575_ (.D(_00429_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[400][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14576_ (.D(_00430_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14577_ (.D(_00431_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14578_ (.D(_00432_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[398][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14579_ (.D(_00433_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[398][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14580_ (.D(_00434_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[397][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14581_ (.D(_00435_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[397][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14582_ (.D(_00436_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[396][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14583_ (.D(_00437_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[396][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14584_ (.D(_00438_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[395][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14585_ (.D(_00439_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[395][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14586_ (.D(_00440_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[394][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14587_ (.D(_00441_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[394][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14588_ (.D(_00442_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[393][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14589_ (.D(_00443_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[393][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14590_ (.D(_00444_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[392][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14591_ (.D(_00445_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[392][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14592_ (.D(_00446_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[391][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14593_ (.D(_00447_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[391][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14594_ (.D(_00448_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[390][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14595_ (.D(_00449_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[390][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14596_ (.D(_00450_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[38][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14597_ (.D(_00451_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[38][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14598_ (.D(_00452_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[388][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14599_ (.D(_00453_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[388][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14600_ (.D(_00454_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[387][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14601_ (.D(_00455_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[387][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14602_ (.D(_00456_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[386][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14603_ (.D(_00457_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[386][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14604_ (.D(_00458_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[385][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14605_ (.D(_00459_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[385][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14606_ (.D(_00460_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[384][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14607_ (.D(_00461_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[384][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14608_ (.D(_00462_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[383][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14609_ (.D(_00463_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[383][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14610_ (.D(_00464_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[382][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14611_ (.D(_00465_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[382][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14612_ (.D(_00466_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[381][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14613_ (.D(_00467_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[381][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14614_ (.D(_00468_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[380][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14615_ (.D(_00469_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[380][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14616_ (.D(_00470_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[37][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14617_ (.D(_00471_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[37][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14618_ (.D(_00472_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[378][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14619_ (.D(_00473_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[378][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14620_ (.D(_00474_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[377][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14621_ (.D(_00475_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[377][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14622_ (.D(_00476_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[376][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14623_ (.D(_00477_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[376][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14624_ (.D(_00478_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[375][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14625_ (.D(_00479_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[375][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14626_ (.D(_00480_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[374][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14627_ (.D(_00481_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[374][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14628_ (.D(_00482_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[373][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14629_ (.D(_00483_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[373][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14630_ (.D(_00484_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[372][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14631_ (.D(_00485_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[372][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14632_ (.D(_00486_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[371][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14633_ (.D(_00487_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[371][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14634_ (.D(_00488_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[370][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14635_ (.D(_00489_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[370][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14636_ (.D(_00490_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[36][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14637_ (.D(_00491_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[36][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14638_ (.D(_00492_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[368][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14639_ (.D(_00493_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[368][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14640_ (.D(_00494_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[367][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14641_ (.D(_00495_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[367][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14642_ (.D(_00496_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[366][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14643_ (.D(_00497_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[366][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14644_ (.D(_00498_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[365][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14645_ (.D(_00499_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[365][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14646_ (.D(_00500_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[364][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14647_ (.D(_00501_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[364][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14648_ (.D(_00502_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[363][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14649_ (.D(_00503_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[363][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14650_ (.D(_00504_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[362][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14651_ (.D(_00505_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[362][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14652_ (.D(_00506_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[361][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14653_ (.D(_00507_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[361][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14654_ (.D(_00508_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[360][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14655_ (.D(_00509_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[360][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14656_ (.D(_00510_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[35][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14657_ (.D(_00511_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[35][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14658_ (.D(_00512_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[358][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14659_ (.D(_00513_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[358][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14660_ (.D(_00514_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[357][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14661_ (.D(_00515_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[357][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14662_ (.D(_00516_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[356][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14663_ (.D(_00517_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[356][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14664_ (.D(_00518_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[355][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14665_ (.D(_00519_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[355][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14666_ (.D(_00520_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[354][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14667_ (.D(_00521_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[354][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14668_ (.D(_00522_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[353][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14669_ (.D(_00523_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[353][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14670_ (.D(_00524_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[352][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14671_ (.D(_00525_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[352][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14672_ (.D(_00526_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[351][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14673_ (.D(_00527_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[351][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14674_ (.D(_00528_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[350][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14675_ (.D(_00529_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[350][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14676_ (.D(_00530_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[34][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14677_ (.D(_00531_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[34][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14678_ (.D(_00532_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[348][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14679_ (.D(_00533_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[348][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14680_ (.D(_00534_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[347][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14681_ (.D(_00535_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[347][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14682_ (.D(_00536_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[346][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14683_ (.D(_00537_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[346][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14684_ (.D(_00538_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[345][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14685_ (.D(_00539_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[345][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14686_ (.D(_00540_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[344][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14687_ (.D(_00541_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[344][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14688_ (.D(_00542_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[343][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14689_ (.D(_00543_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[343][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14690_ (.D(_00544_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[342][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14691_ (.D(_00545_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[342][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14692_ (.D(_00546_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[341][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14693_ (.D(_00547_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[341][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14694_ (.D(_00548_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[340][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14695_ (.D(_00549_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[340][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14696_ (.D(_00550_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[33][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14697_ (.D(_00551_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[33][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14698_ (.D(_00552_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[338][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14699_ (.D(_00553_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[338][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14700_ (.D(_00554_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[337][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14701_ (.D(_00555_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[337][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14702_ (.D(_00556_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[336][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14703_ (.D(_00557_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[336][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14704_ (.D(_00558_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[335][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14705_ (.D(_00559_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[335][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14706_ (.D(_00560_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[334][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14707_ (.D(_00561_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[334][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14708_ (.D(_00562_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[333][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14709_ (.D(_00563_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[333][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14710_ (.D(_00564_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[332][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14711_ (.D(_00565_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[332][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14712_ (.D(_00566_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[331][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14713_ (.D(_00567_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[331][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14714_ (.D(_00568_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[330][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14715_ (.D(_00569_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[330][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14716_ (.D(_00570_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[32][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14717_ (.D(_00571_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[32][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14718_ (.D(_00572_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[328][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14719_ (.D(_00573_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[328][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14720_ (.D(_00574_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[327][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14721_ (.D(_00575_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[327][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14722_ (.D(_00576_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[326][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14723_ (.D(_00577_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[326][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14724_ (.D(_00578_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[325][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14725_ (.D(_00579_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[325][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14726_ (.D(_00580_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[324][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14727_ (.D(_00581_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[324][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14728_ (.D(_00582_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[323][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14729_ (.D(_00583_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[323][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14730_ (.D(_00584_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[322][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14731_ (.D(_00585_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[322][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14732_ (.D(_00586_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[321][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14733_ (.D(_00587_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[321][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14734_ (.D(_00588_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[320][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14735_ (.D(_00589_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[320][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14736_ (.D(_00590_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[31][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14737_ (.D(_00591_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[31][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14738_ (.D(_00592_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[318][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14739_ (.D(_00593_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[318][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14740_ (.D(_00594_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[317][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14741_ (.D(_00595_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[317][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14742_ (.D(_00596_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[316][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14743_ (.D(_00597_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[316][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14744_ (.D(_00598_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[315][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14745_ (.D(_00599_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[315][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14746_ (.D(_00600_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[314][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14747_ (.D(_00601_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[314][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14748_ (.D(_00602_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[313][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14749_ (.D(_00603_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[313][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14750_ (.D(_00604_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[312][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14751_ (.D(_00605_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[312][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14752_ (.D(_00606_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[311][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14753_ (.D(_00607_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[311][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14754_ (.D(_00608_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[310][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14755_ (.D(_00609_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[310][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14756_ (.D(_00610_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[30][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14757_ (.D(_00611_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[30][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14758_ (.D(_00612_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[308][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14759_ (.D(_00613_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[308][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14760_ (.D(_00614_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[307][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14761_ (.D(_00615_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[307][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14762_ (.D(_00616_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[306][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14763_ (.D(_00617_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[306][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14764_ (.D(_00618_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[305][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14765_ (.D(_00619_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[305][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14766_ (.D(_00620_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[304][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14767_ (.D(_00621_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[304][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14768_ (.D(_00622_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[303][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14769_ (.D(_00623_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[303][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14770_ (.D(_00624_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[302][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14771_ (.D(_00625_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[302][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14772_ (.D(_00626_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[301][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14773_ (.D(_00627_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[301][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14774_ (.D(_00628_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[300][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14775_ (.D(_00629_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[300][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14776_ (.D(_00630_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14777_ (.D(_00631_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14778_ (.D(_00632_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[298][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14779_ (.D(_00633_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[298][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14780_ (.D(_00634_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[297][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14781_ (.D(_00635_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[297][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14782_ (.D(_00636_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[296][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14783_ (.D(_00637_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[296][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14784_ (.D(_00638_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[295][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14785_ (.D(_00639_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[295][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14786_ (.D(_00640_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[294][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14787_ (.D(_00641_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[294][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14788_ (.D(_00642_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[293][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14789_ (.D(_00643_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[293][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14790_ (.D(_00644_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[292][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14791_ (.D(_00645_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[292][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14792_ (.D(_00646_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[291][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14793_ (.D(_00647_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[291][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14794_ (.D(_00648_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[290][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14795_ (.D(_00649_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[290][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14796_ (.D(_00650_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[28][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14797_ (.D(_00651_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[28][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14798_ (.D(_00652_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[288][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14799_ (.D(_00653_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[288][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14800_ (.D(_00654_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[287][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14801_ (.D(_00655_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[287][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14802_ (.D(_00656_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[286][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14803_ (.D(_00657_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[286][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14804_ (.D(_00658_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[285][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14805_ (.D(_00659_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[285][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14806_ (.D(_00660_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[284][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14807_ (.D(_00661_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[284][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14808_ (.D(_00662_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[283][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14809_ (.D(_00663_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[283][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14810_ (.D(_00664_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[282][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14811_ (.D(_00665_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[282][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14812_ (.D(_00666_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[281][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14813_ (.D(_00667_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[281][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14814_ (.D(_00668_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[280][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14815_ (.D(_00669_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[280][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14816_ (.D(_00670_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[27][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14817_ (.D(_00671_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[27][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14818_ (.D(_00672_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[278][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14819_ (.D(_00673_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[278][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14820_ (.D(_00674_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[277][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14821_ (.D(_00675_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[277][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14822_ (.D(_00676_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[276][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14823_ (.D(_00677_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[276][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14824_ (.D(_00678_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[275][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14825_ (.D(_00679_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[275][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14826_ (.D(_00680_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[274][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14827_ (.D(_00681_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[274][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14828_ (.D(_00682_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[273][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14829_ (.D(_00683_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[273][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14830_ (.D(_00684_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[272][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14831_ (.D(_00685_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[272][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14832_ (.D(_00686_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[271][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14833_ (.D(_00687_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[271][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14834_ (.D(_00688_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[270][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14835_ (.D(_00689_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[270][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14836_ (.D(_00690_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[26][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14837_ (.D(_00691_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[26][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14838_ (.D(_00692_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[268][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14839_ (.D(_00693_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[268][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14840_ (.D(_00694_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[267][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14841_ (.D(_00695_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[267][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14842_ (.D(_00696_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[266][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14843_ (.D(_00697_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[266][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14844_ (.D(_00698_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[265][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14845_ (.D(_00699_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[265][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14846_ (.D(_00700_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[264][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14847_ (.D(_00701_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[264][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14848_ (.D(_00702_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[263][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14849_ (.D(_00703_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[263][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14850_ (.D(_00704_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[262][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14851_ (.D(_00705_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[262][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14852_ (.D(_00706_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[261][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14853_ (.D(_00707_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[261][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14854_ (.D(_00708_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[260][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14855_ (.D(_00709_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[260][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14856_ (.D(_00710_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[25][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14857_ (.D(_00711_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[25][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14858_ (.D(_00712_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[24][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14859_ (.D(_00713_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[24][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14860_ (.D(_00714_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[258][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14861_ (.D(_00715_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[258][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14862_ (.D(_00716_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[257][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14863_ (.D(_00717_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[257][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14864_ (.D(_00718_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[250][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14865_ (.D(_00719_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[250][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14866_ (.D(_00720_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[256][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14867_ (.D(_00721_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[256][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14868_ (.D(_00722_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[255][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14869_ (.D(_00723_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[255][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14870_ (.D(_00724_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[251][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14871_ (.D(_00725_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[251][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14872_ (.D(_00726_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[254][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14873_ (.D(_00727_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[254][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14874_ (.D(_00728_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[252][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14875_ (.D(_00729_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[252][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14876_ (.D(_00730_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[253][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14877_ (.D(_00731_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[253][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14878_ (.D(_00732_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[248][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14879_ (.D(_00733_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[248][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14880_ (.D(_00734_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[243][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14881_ (.D(_00735_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[243][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14882_ (.D(_00736_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[242][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14883_ (.D(_00737_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[242][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14884_ (.D(_00738_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[241][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14885_ (.D(_00739_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[241][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14886_ (.D(_00740_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[240][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14887_ (.D(_00741_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[240][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14888_ (.D(_00742_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[23][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14889_ (.D(_00743_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[23][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14890_ (.D(_00744_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[238][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14891_ (.D(_00745_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[238][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14892_ (.D(_00746_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[239][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14893_ (.D(_00747_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[239][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14894_ (.D(_00748_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[237][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14895_ (.D(_00749_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[237][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14896_ (.D(_00750_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[236][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14897_ (.D(_00751_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[236][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14898_ (.D(_00752_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[235][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14899_ (.D(_00753_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[235][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14900_ (.D(_00754_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[234][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14901_ (.D(_00755_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[234][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14902_ (.D(_00756_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[233][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14903_ (.D(_00757_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[233][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14904_ (.D(_00758_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[232][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14905_ (.D(_00759_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[232][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14906_ (.D(_00760_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[231][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14907_ (.D(_00761_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[231][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14908_ (.D(_00762_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[49][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14909_ (.D(_00763_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[49][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14910_ (.D(_00764_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[230][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14911_ (.D(_00765_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[230][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14912_ (.D(_00766_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[22][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14913_ (.D(_00767_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[22][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14914_ (.D(_00768_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[39][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14915_ (.D(_00769_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[39][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14916_ (.D(_00770_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[228][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14917_ (.D(_00771_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[228][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14918_ (.D(_00772_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[159][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14919_ (.D(_00773_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[159][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14920_ (.D(_00774_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[149][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14921_ (.D(_00775_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[149][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14922_ (.D(_00776_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14923_ (.D(_00777_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14924_ (.D(_00778_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[70][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14925_ (.D(_00779_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[70][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14926_ (.D(_00780_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[72][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14927_ (.D(_00781_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[72][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14928_ (.D(_00782_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[71][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14929_ (.D(_00783_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[71][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14930_ (.D(_00784_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[227][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14931_ (.D(_00785_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[227][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14932_ (.D(_00786_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[226][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14933_ (.D(_00787_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[226][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14934_ (.D(_00788_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[225][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14935_ (.D(_00789_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[225][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14936_ (.D(_00790_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[224][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14937_ (.D(_00791_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[224][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14938_ (.D(_00792_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[223][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14939_ (.D(_00793_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[223][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14940_ (.D(_00794_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[222][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14941_ (.D(_00795_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[222][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14942_ (.D(_00796_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[221][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14943_ (.D(_00797_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[221][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14944_ (.D(_00798_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[169][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14945_ (.D(_00799_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[169][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14946_ (.D(_00800_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[220][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14947_ (.D(_00801_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[220][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14948_ (.D(_00802_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[21][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14949_ (.D(_00803_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[21][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14950_ (.D(_00804_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[218][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14951_ (.D(_00805_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[218][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14952_ (.D(_00806_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[529][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14953_ (.D(_00807_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[529][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14954_ (.D(_00808_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[539][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14955_ (.D(_00809_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[539][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14956_ (.D(_00810_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[217][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14957_ (.D(_00811_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[217][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14958_ (.D(_00812_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[549][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14959_ (.D(_00813_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[549][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14960_ (.D(_00814_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[216][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14961_ (.D(_00815_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[216][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14962_ (.D(_00816_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[559][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14963_ (.D(_00817_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[559][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14964_ (.D(_00818_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[569][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14965_ (.D(_00819_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[569][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14966_ (.D(_00820_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[215][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14967_ (.D(_00821_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[215][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14968_ (.D(_00822_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[575][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14969_ (.D(_00823_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[575][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14970_ (.D(_00824_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[57][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14971_ (.D(_00825_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[57][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14972_ (.D(_00826_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[214][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14973_ (.D(_00827_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[214][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14974_ (.D(_00828_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[58][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14975_ (.D(_00829_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[58][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14976_ (.D(_00830_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[19][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14977_ (.D(_00831_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[19][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14978_ (.D(_00832_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14979_ (.D(_00833_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14980_ (.D(_00834_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[60][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14981_ (.D(_00835_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[60][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14982_ (.D(_00836_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[213][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14983_ (.D(_00837_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[213][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14984_ (.D(_00838_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[61][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14985_ (.D(_00839_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[61][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14986_ (.D(_00840_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[62][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14987_ (.D(_00841_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[62][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14988_ (.D(_00842_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[29][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14989_ (.D(_00843_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[29][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14990_ (.D(_00844_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[63][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14991_ (.D(_00845_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[63][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14992_ (.D(_00846_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[64][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14993_ (.D(_00847_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[64][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14994_ (.D(_00848_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[212][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14995_ (.D(_00849_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[212][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14996_ (.D(_00850_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[65][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14997_ (.D(_00851_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[65][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14998_ (.D(_00852_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[66][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _14999_ (.D(_00853_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[66][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15000_ (.D(_00854_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[67][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15001_ (.D(_00855_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[67][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15002_ (.D(_00856_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[211][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15003_ (.D(_00857_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[211][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15004_ (.D(_00858_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[68][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15005_ (.D(_00859_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[68][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15006_ (.D(_00860_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[210][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15007_ (.D(_00861_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[210][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15008_ (.D(_00862_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[20][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15009_ (.D(_00863_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[20][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15010_ (.D(_00864_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[208][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15011_ (.D(_00865_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[208][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15012_ (.D(_00866_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[74][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15013_ (.D(_00867_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[74][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15014_ (.D(_00868_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[75][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15015_ (.D(_00869_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[75][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15016_ (.D(_00870_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[207][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15017_ (.D(_00871_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[207][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15018_ (.D(_00872_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[206][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15019_ (.D(_00873_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[206][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15020_ (.D(_00874_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[73][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15021_ (.D(_00875_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[73][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15022_ (.D(_00876_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[205][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15023_ (.D(_00877_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[205][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15024_ (.D(_00878_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[76][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15025_ (.D(_00879_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[76][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15026_ (.D(_00880_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[204][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15027_ (.D(_00881_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[204][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15028_ (.D(_00882_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[203][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15029_ (.D(_00883_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[203][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15030_ (.D(_00884_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[202][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15031_ (.D(_00885_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[202][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15032_ (.D(_00886_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[201][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15033_ (.D(_00887_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[201][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15034_ (.D(_00888_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[200][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15035_ (.D(_00889_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[200][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15036_ (.D(_00890_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15037_ (.D(_00891_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15038_ (.D(_00892_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[198][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15039_ (.D(_00893_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[198][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15040_ (.D(_00894_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[119][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15041_ (.D(_00895_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[119][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15042_ (.D(_00896_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[197][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15043_ (.D(_00897_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[197][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15044_ (.D(_00898_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[109][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15045_ (.D(_00899_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[109][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15046_ (.D(_00900_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[196][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15047_ (.D(_00901_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[196][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15048_ (.D(_00902_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[195][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15049_ (.D(_00903_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[195][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15050_ (.D(_00904_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[194][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15051_ (.D(_00905_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[194][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15052_ (.D(_00906_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[193][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15053_ (.D(_00907_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[193][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15054_ (.D(_00908_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[192][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15055_ (.D(_00909_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[192][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15056_ (.D(_00910_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[191][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15057_ (.D(_00911_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[191][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15058_ (.D(_00912_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[190][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15059_ (.D(_00913_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[190][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15060_ (.D(_00914_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[18][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15061_ (.D(_00915_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[18][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15062_ (.D(_00916_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[188][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15063_ (.D(_00917_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[188][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15064_ (.D(_00918_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[187][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15065_ (.D(_00919_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[187][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15066_ (.D(_00920_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[186][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15067_ (.D(_00921_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[186][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15068_ (.D(_00922_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[185][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15069_ (.D(_00923_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[185][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15070_ (.D(_00924_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[189][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15071_ (.D(_00925_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[189][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15072_ (.D(_00926_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[179][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15073_ (.D(_00927_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[179][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15074_ (.D(_00928_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[184][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15075_ (.D(_00929_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[184][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15076_ (.D(_00930_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[183][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15077_ (.D(_00931_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[183][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15078_ (.D(_00932_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[182][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15079_ (.D(_00933_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[182][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15080_ (.D(_00934_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[181][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15081_ (.D(_00935_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[181][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15082_ (.D(_00936_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[122][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15083_ (.D(_00937_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[122][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15084_ (.D(_00938_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[180][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15085_ (.D(_00939_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[180][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15086_ (.D(_00940_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[499][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15087_ (.D(_00941_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[499][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15088_ (.D(_00942_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[17][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15089_ (.D(_00943_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[17][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15090_ (.D(_00944_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[178][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15091_ (.D(_00945_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[178][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15092_ (.D(_00946_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[177][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15093_ (.D(_00947_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[177][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15094_ (.D(_00948_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[509][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15095_ (.D(_00949_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[509][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15096_ (.D(_00950_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[479][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15097_ (.D(_00951_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[479][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15098_ (.D(_00952_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[176][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15099_ (.D(_00953_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[176][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15100_ (.D(_00954_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[175][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15101_ (.D(_00955_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[175][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15102_ (.D(_00956_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[489][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15103_ (.D(_00957_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[489][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15104_ (.D(_00958_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[174][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15105_ (.D(_00959_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[174][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15106_ (.D(_00960_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[439][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15107_ (.D(_00961_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[439][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15108_ (.D(_00962_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[173][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15109_ (.D(_00963_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[173][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15110_ (.D(_00964_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[172][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15111_ (.D(_00965_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[172][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15112_ (.D(_00966_),
    .CLK(net3),
    .Q(\mod.u_cpu.raddr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15113_ (.D(_00002_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15114_ (.D(_00967_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[419][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15115_ (.D(_00968_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[419][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15116_ (.D(_00969_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[519][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15117_ (.D(_00970_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[519][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15118_ (.D(_00971_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[449][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15119_ (.D(_00972_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[449][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15120_ (.D(_00973_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[171][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15121_ (.D(_00974_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[171][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15122_ (.D(_00975_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[170][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15123_ (.D(_00976_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[170][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15124_ (.D(_00977_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[459][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15125_ (.D(_00978_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[459][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15126_ (.D(_00979_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[16][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15127_ (.D(_00980_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[16][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15128_ (.D(_00981_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[168][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15129_ (.D(_00982_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[168][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15130_ (.D(_00983_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[167][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15131_ (.D(_00984_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[167][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15132_ (.D(_00985_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[166][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15133_ (.D(_00986_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[166][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15134_ (.D(_00987_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[469][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15135_ (.D(_00988_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[469][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15136_ (.D(_00989_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[429][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15137_ (.D(_00990_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[429][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15138_ (.D(_00991_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[165][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15139_ (.D(_00992_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[165][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15140_ (.D(_00993_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[164][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15141_ (.D(_00994_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[164][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15142_ (.D(_00995_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[163][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15143_ (.D(_00996_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[163][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15144_ (.D(_00997_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[162][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15145_ (.D(_00998_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[162][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15146_ (.D(_00999_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[161][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15147_ (.D(_01000_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[161][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15148_ (.D(_01001_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[160][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15149_ (.D(_01002_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[160][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15150_ (.D(_01003_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15151_ (.D(_01004_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15152_ (.D(_01005_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[158][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15153_ (.D(_01006_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[158][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15154_ (.D(_01007_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[157][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15155_ (.D(_01008_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[157][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15156_ (.D(_01009_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[156][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15157_ (.D(_01010_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[156][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15158_ (.D(_01011_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[155][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15159_ (.D(_01012_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[155][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15160_ (.D(_01013_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[154][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15161_ (.D(_01014_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[154][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15162_ (.D(_01015_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[153][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15163_ (.D(_01016_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[153][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15164_ (.D(_01017_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[152][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15165_ (.D(_01018_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[152][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15166_ (.D(_01019_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[151][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15167_ (.D(_01020_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[151][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15168_ (.D(_01021_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[150][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15169_ (.D(_01022_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[150][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15170_ (.D(_01023_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15171_ (.D(_01024_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15172_ (.D(_01025_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[148][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15173_ (.D(_01026_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[148][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15174_ (.D(_01027_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[147][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15175_ (.D(_01028_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[147][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15176_ (.D(_01029_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[146][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15177_ (.D(_01030_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[146][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15178_ (.D(_01031_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[145][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15179_ (.D(_01032_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[145][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15180_ (.D(_01033_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[144][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15181_ (.D(_01034_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[144][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15182_ (.D(_01035_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[121][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15183_ (.D(_01036_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[121][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15184_ (.D(_01037_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[143][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15185_ (.D(_01038_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[143][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15186_ (.D(_01039_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[142][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15187_ (.D(_01040_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[142][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15188_ (.D(_01041_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[77][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15189_ (.D(_01042_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[77][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15190_ (.D(_01043_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[141][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15191_ (.D(_01044_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[141][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15192_ (.D(_01045_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[140][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15193_ (.D(_01046_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[140][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15194_ (.D(_01047_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15195_ (.D(_01048_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15196_ (.D(_01049_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15197_ (.D(_01050_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15198_ (.D(_01051_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[138][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15199_ (.D(_01052_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[138][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15200_ (.D(_01053_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[137][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15201_ (.D(_01054_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[137][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15202_ (.D(_01055_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[78][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15203_ (.D(_01056_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[78][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15204_ (.D(_01057_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[136][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15205_ (.D(_01058_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[136][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15206_ (.D(_01059_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[209][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15207_ (.D(_01060_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[209][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15208_ (.D(_01061_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[219][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15209_ (.D(_01062_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[219][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15210_ (.D(_01063_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[199][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15211_ (.D(_01064_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[199][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15212_ (.D(_01065_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[80][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15213_ (.D(_01066_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[80][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15214_ (.D(_01067_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[135][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15215_ (.D(_01068_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[135][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15216_ (.D(_01069_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[134][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15217_ (.D(_01070_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[134][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15218_ (.D(_01071_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[133][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15219_ (.D(_01072_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[133][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15220_ (.D(_01073_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[132][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15221_ (.D(_01074_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[132][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15222_ (.D(_01075_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[131][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15223_ (.D(_01076_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[131][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15224_ (.D(_01077_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[130][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15225_ (.D(_01078_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[130][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15226_ (.D(_01079_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15227_ (.D(_01080_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15228_ (.D(_01081_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[128][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15229_ (.D(_01082_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[128][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15230_ (.D(_01083_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[229][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15231_ (.D(_01084_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[229][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15232_ (.D(_01085_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[127][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15233_ (.D(_01086_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[127][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15234_ (.D(_01087_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[126][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15235_ (.D(_01088_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[126][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15236_ (.D(_01089_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[125][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15237_ (.D(_01090_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[125][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15238_ (.D(_01091_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[124][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15239_ (.D(_01092_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[124][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15240_ (.D(_01093_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram_if.rreq_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15241_ (.D(_01094_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[123][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15242_ (.D(_01095_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[123][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15243_ (.D(_00008_),
    .CLK(net4),
    .Q(\mod.timer_irq ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15244_ (.D(_00019_),
    .CLK(net4),
    .Q(\mod.u_arbiter.i_wb_cpu_ack ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15245_ (.D(_00030_),
    .CLK(net4),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15246_ (.D(_00041_),
    .CLK(net4),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15247_ (.D(_00052_),
    .CLK(net4),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15248_ (.D(_00063_),
    .CLK(net4),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15249_ (.D(_00074_),
    .CLK(net4),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15250_ (.D(_00075_),
    .CLK(net4),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15251_ (.D(_00076_),
    .CLK(net4),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15252_ (.D(_00077_),
    .CLK(net4),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15253_ (.D(_00009_),
    .CLK(net4),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15254_ (.D(_00010_),
    .CLK(net4),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15255_ (.D(_00011_),
    .CLK(net4),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15256_ (.D(_00012_),
    .CLK(net4),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15257_ (.D(_00013_),
    .CLK(net4),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15258_ (.D(_00014_),
    .CLK(net4),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15259_ (.D(_00015_),
    .CLK(net4),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15260_ (.D(_00016_),
    .CLK(net4),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15261_ (.D(_00017_),
    .CLK(net4),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15262_ (.D(_00018_),
    .CLK(net4),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15263_ (.D(_00020_),
    .CLK(net4),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15264_ (.D(_00021_),
    .CLK(net4),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15265_ (.D(_00022_),
    .CLK(net4),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15266_ (.D(_00023_),
    .CLK(net4),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15267_ (.D(_00024_),
    .CLK(net4),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15268_ (.D(_00025_),
    .CLK(net4),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15269_ (.D(_00026_),
    .CLK(net4),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15270_ (.D(_00027_),
    .CLK(net4),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15271_ (.D(_00028_),
    .CLK(net4),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15272_ (.D(_00029_),
    .CLK(net4),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15273_ (.D(_00031_),
    .CLK(net4),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15274_ (.D(_00032_),
    .CLK(net4),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15275_ (.D(_00033_),
    .CLK(net4),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15276_ (.D(_00034_),
    .CLK(net4),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15277_ (.D(_00035_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[34] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15278_ (.D(_00036_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[35] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15279_ (.D(_00037_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[36] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15280_ (.D(_00038_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[37] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15281_ (.D(_00039_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[38] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15282_ (.D(_00040_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[39] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15283_ (.D(_00042_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[40] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15284_ (.D(_00043_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[41] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15285_ (.D(_00044_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[42] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15286_ (.D(_00045_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[43] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15287_ (.D(_00046_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[44] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15288_ (.D(_00047_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[45] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15289_ (.D(_00048_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[46] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15290_ (.D(_00049_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[47] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15291_ (.D(_00050_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[48] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15292_ (.D(_00051_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[49] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15293_ (.D(_00053_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[50] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15294_ (.D(_00054_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[51] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15295_ (.D(_00055_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[52] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15296_ (.D(_00056_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[53] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15297_ (.D(_00057_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[54] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15298_ (.D(_00058_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[55] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15299_ (.D(_00059_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[56] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15300_ (.D(_00060_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[57] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15301_ (.D(_00061_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[58] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15302_ (.D(_00062_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[59] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15303_ (.D(_00064_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[60] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15304_ (.D(_00065_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[61] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15305_ (.D(_00066_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[62] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15306_ (.D(_00067_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[63] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15307_ (.D(_00068_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[64] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15308_ (.D(_00069_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[65] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15309_ (.D(_00070_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[66] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15310_ (.D(_00071_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[67] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15311_ (.D(_00072_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[68] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15312_ (.D(_00073_),
    .CLK(net4),
    .Q(\mod.u_scanchain_local.module_data_in[69] ));
 gf180mcu_fd_sc_mcu7t5v0__dffnq_1 _15313_ (.D(\mod.u_scanchain_local.module_data_in[69] ),
    .CLKN(net4),
    .Q(net7));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15314_ (.D(\mod.u_cpu.cpu.o_wen0 ),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram_if.wen0_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15315_ (.D(\mod.u_cpu.rf_ram_if.wdata1_r[1] ),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram_if.wdata1_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15316_ (.D(\mod.u_cpu.cpu.o_wdata1 ),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram_if.wdata1_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15317_ (.D(_01096_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15318_ (.D(_01097_),
    .CLK(net3),
    .Q(\mod.u_cpu.raddr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15319_ (.D(_01098_),
    .CLK(net3),
    .Q(\mod.u_cpu.raddr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15320_ (.D(_01099_),
    .CLK(net3),
    .Q(\mod.u_cpu.raddr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15321_ (.D(\mod.u_cpu.rf_ram_if.rtrig0 ),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram_if.rtrig1 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15322_ (.D(_01100_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram_if.rgnt ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15323_ (.D(_01101_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram_if.rdata0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15324_ (.D(_01102_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram_if.rdata1 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15325_ (.D(\mod.u_cpu.cpu.o_wdata0 ),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram_if.wdata0_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15326_ (.D(_01103_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.state.ibus_cyc ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15327_ (.D(_01104_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[409][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15328_ (.D(_01105_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[409][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15329_ (.D(\mod.u_cpu.cpu.o_wen1 ),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram_if.wen1_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15330_ (.D(_01106_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[246][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15331_ (.D(_01107_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[246][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15332_ (.D(_00007_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.regzero ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15333_ (.D(_01108_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[99][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15334_ (.D(_01109_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[99][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15335_ (.D(_01110_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[89][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15336_ (.D(_01111_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[89][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15337_ (.D(_01112_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[98][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15338_ (.D(_01113_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[98][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15339_ (.D(_01114_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[96][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15340_ (.D(_01115_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[96][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15341_ (.D(_01116_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[97][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15342_ (.D(_01117_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[97][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15343_ (.D(_01118_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[399][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15344_ (.D(_01119_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[399][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15345_ (.D(_01120_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[389][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15346_ (.D(_01121_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[389][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15347_ (.D(_01122_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[379][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15348_ (.D(_01123_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[379][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15349_ (.D(_01124_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[369][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15350_ (.D(_01125_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[369][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15351_ (.D(_01126_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.genblk3.csr.o_new_irq ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15352_ (.D(_01127_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.ctrl.i_iscomp ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15353_ (.D(_01128_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.genblk3.csr.mstatus_mie ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15354_ (.D(_01129_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.genblk3.csr.mie_mtie ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15355_ (.D(_01130_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.genblk3.csr.mstatus_mpie ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15356_ (.D(_01131_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.genblk3.csr.mcause31 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15357_ (.D(_01132_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.genblk3.csr.mcause3_0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15358_ (.D(_01133_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.genblk3.csr.mcause3_0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15359_ (.D(_01134_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.genblk3.csr.mcause3_0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15360_ (.D(_01135_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.genblk3.csr.mcause3_0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15361_ (.D(_01136_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[86][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15362_ (.D(_01137_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[86][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15363_ (.D(_01138_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[85][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15364_ (.D(_01139_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[85][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15365_ (.D(_01140_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15366_ (.D(_01141_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[10][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15367_ (.D(_01142_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[84][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15368_ (.D(_01143_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[84][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15369_ (.D(_01144_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[108][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15370_ (.D(_01145_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[108][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15371_ (.D(_01146_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[83][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15372_ (.D(_01147_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[83][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15373_ (.D(_01148_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[107][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15374_ (.D(_01149_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[107][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15375_ (.D(_01150_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[79][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15376_ (.D(_01151_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[79][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15377_ (.D(_01152_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[82][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15378_ (.D(_01153_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[82][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15379_ (.D(_01154_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[69][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15380_ (.D(_01155_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[69][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15381_ (.D(_01156_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[106][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15382_ (.D(_01157_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[106][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15383_ (.D(_01158_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[81][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15384_ (.D(_01159_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[81][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15385_ (.D(_01160_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[105][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15386_ (.D(_01161_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[105][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15387_ (.D(_01162_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[104][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15388_ (.D(_01163_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[104][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15389_ (.D(_01164_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[103][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15390_ (.D(_01165_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[103][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15391_ (.D(_01166_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[59][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15392_ (.D(_01167_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[59][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15393_ (.D(_01168_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[102][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15394_ (.D(_01169_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[102][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15395_ (.D(_01170_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[101][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15396_ (.D(_01171_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[101][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15397_ (.D(_01172_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[100][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15398_ (.D(_01173_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[100][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15399_ (.D(_01174_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15400_ (.D(_01175_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15401_ (.D(_01176_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[359][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15402_ (.D(_01177_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[359][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15403_ (.D(_01178_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15404_ (.D(_01179_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15405_ (.D(_01180_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15406_ (.D(_01181_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15407_ (.D(_01182_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15408_ (.D(_01183_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15409_ (.D(_01184_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15410_ (.D(_01185_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15411_ (.D(_01186_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15412_ (.D(_01187_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15413_ (.D(_01188_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15414_ (.D(_01189_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15415_ (.D(_01190_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15416_ (.D(_01191_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15417_ (.D(_01192_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15418_ (.D(_01193_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15419_ (.D(_01194_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[349][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15420_ (.D(_01195_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[349][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15421_ (.D(_01196_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.genblk1.align.ctrl_misal ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15422_ (.D(_01197_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.bufreg.i_sh_signed ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15423_ (.D(_01198_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[94][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15424_ (.D(_01199_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[94][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15425_ (.D(_01200_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[93][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15426_ (.D(_01201_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[93][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15427_ (.D(_01202_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[92][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15428_ (.D(_01203_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[92][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15429_ (.D(_01204_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[95][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15430_ (.D(_01205_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[95][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15431_ (.D(_01206_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.immdec.imm11_7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15432_ (.D(_01207_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.immdec.imm11_7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15433_ (.D(_01208_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.immdec.imm11_7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15434_ (.D(_01209_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.immdec.imm11_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15435_ (.D(_01210_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.immdec.imm11_7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15436_ (.D(_01211_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[91][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15437_ (.D(_01212_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[91][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15438_ (.D(_01213_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[139][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15439_ (.D(_01214_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[139][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15440_ (.D(_00003_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.alu.add_cy_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15441_ (.D(_01215_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[339][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15442_ (.D(_01216_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[339][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15443_ (.D(_01217_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15444_ (.D(_01218_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15445_ (.D(_01219_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15446_ (.D(_01220_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15447_ (.D(_01221_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15448_ (.D(_01222_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15449_ (.D(_01223_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15450_ (.D(_01224_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15451_ (.D(_01225_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15452_ (.D(_01226_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15453_ (.D(_01227_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15454_ (.D(_01228_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15455_ (.D(_01229_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15456_ (.D(_01230_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15457_ (.D(_01231_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15458_ (.D(_01232_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15459_ (.D(_01233_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15460_ (.D(_01234_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15461_ (.D(_01235_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15462_ (.D(_01236_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15463_ (.D(_01237_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15464_ (.D(_01238_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15465_ (.D(_01239_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15466_ (.D(_01240_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15467_ (.D(_01241_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15468_ (.D(_01242_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15469_ (.D(_01243_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15470_ (.D(_01244_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15471_ (.D(_01245_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15472_ (.D(_01246_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15473_ (.D(_01247_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15474_ (.D(_01248_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15475_ (.D(_00005_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.ctrl.pc_plus_4_cy_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15476_ (.D(_00006_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.ctrl.pc_plus_offset_cy_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15477_ (.D(_01249_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.bufreg.lsb[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15478_ (.D(_01250_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.bufreg.lsb[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15479_ (.D(_01251_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[129][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15480_ (.D(_01252_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[129][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15481_ (.D(_00004_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.bufreg.c_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15482_ (.D(_01253_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15483_ (.D(_01254_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15484_ (.D(_01255_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15485_ (.D(_01256_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15486_ (.D(_01257_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15487_ (.D(_01258_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15488_ (.D(_01259_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15489_ (.D(_01260_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15490_ (.D(_01261_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15491_ (.D(_01262_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15492_ (.D(_01263_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15493_ (.D(_01264_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15494_ (.D(_01265_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15495_ (.D(_01266_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15496_ (.D(_01267_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15497_ (.D(_01268_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15498_ (.D(_01269_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15499_ (.D(_01270_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15500_ (.D(_01271_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15501_ (.D(_01272_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15502_ (.D(_01273_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15503_ (.D(_01274_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15504_ (.D(_01275_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15505_ (.D(_01276_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15506_ (.D(_01277_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15507_ (.D(_01278_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15508_ (.D(_01279_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15509_ (.D(_01280_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15510_ (.D(_01281_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15511_ (.D(_01282_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15512_ (.D(_01283_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[329][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15513_ (.D(_01284_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[329][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15514_ (.D(_01285_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.alu.cmp_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15515_ (.D(_01286_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[319][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15516_ (.D(_01287_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[319][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15517_ (.D(_01288_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[309][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15518_ (.D(_01289_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[309][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15519_ (.D(_01290_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.genblk3.csr.timer_irq_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15520_ (.D(_01291_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.immdec.imm31 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15521_ (.D(_01292_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.immdec.imm19_12_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15522_ (.D(_01293_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.immdec.imm19_12_20[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15523_ (.D(_01294_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.immdec.imm19_12_20[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15524_ (.D(_01295_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.immdec.imm19_12_20[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15525_ (.D(_01296_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.csr_imm ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15526_ (.D(_01297_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.immdec.imm19_12_20[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15527_ (.D(_01298_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.immdec.imm19_12_20[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15528_ (.D(_01299_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.immdec.imm19_12_20[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15529_ (.D(_01300_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.immdec.imm19_12_20[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15530_ (.D(_01301_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.immdec.imm7 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15531_ (.D(_01302_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.immdec.imm30_25[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15532_ (.D(_01303_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.immdec.imm30_25[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15533_ (.D(_01304_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.immdec.imm30_25[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15534_ (.D(_01305_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.immdec.imm30_25[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15535_ (.D(_01306_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.immdec.imm30_25[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15536_ (.D(_01307_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.immdec.imm30_25[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15537_ (.D(_01308_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15538_ (.D(_01309_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.immdec.imm24_20[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15539_ (.D(_01310_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.immdec.imm24_20[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15540_ (.D(_01311_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.immdec.imm24_20[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15541_ (.D(_01312_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.immdec.imm24_20[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15542_ (.D(_01313_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.decode.op26 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15543_ (.D(_01314_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[112][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15544_ (.D(_01315_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[112][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15545_ (.D(_01316_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.decode.op22 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15546_ (.D(_01317_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.decode.op21 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15547_ (.D(_01318_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15548_ (.D(_01319_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15549_ (.D(_01320_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.decode.co_mem_word ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15550_ (.D(_01321_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.csr_d_sel ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15551_ (.D(_01322_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.decode.opcode[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15552_ (.D(_01323_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.decode.opcode[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15553_ (.D(_01324_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.decode.opcode[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15554_ (.D(_01325_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_we ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15555_ (.D(_01326_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.branch_op ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15556_ (.D(_01327_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[111][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15557_ (.D(_01328_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[111][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15558_ (.D(_01329_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15559_ (.D(_01330_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15560_ (.D(_01331_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15561_ (.D(_01332_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15562_ (.D(_01333_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15563_ (.D(_01334_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15564_ (.D(_01335_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15565_ (.D(_01336_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15566_ (.D(_01337_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15567_ (.D(_01338_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15568_ (.D(_01339_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15569_ (.D(_01340_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15570_ (.D(_01341_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15571_ (.D(_01342_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15572_ (.D(_01343_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15573_ (.D(_01344_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15574_ (.D(_01345_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15575_ (.D(_01346_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15576_ (.D(_01347_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15577_ (.D(_01348_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15578_ (.D(_01349_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15579_ (.D(_01350_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15580_ (.D(_01351_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15581_ (.D(_01352_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15582_ (.D(_01353_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15583_ (.D(_01354_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15584_ (.D(_01355_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15585_ (.D(_01356_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15586_ (.D(_01357_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15587_ (.D(_01358_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15588_ (.D(_01359_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15589_ (.D(_01360_),
    .CLK(net3),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15590_ (.D(_01361_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[114][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15591_ (.D(_01362_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[114][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15592_ (.D(_01363_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[299][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15593_ (.D(_01364_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[299][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15594_ (.D(_01365_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[113][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15595_ (.D(_01366_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[113][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15596_ (.D(_01367_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[245][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15597_ (.D(_01368_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[245][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15598_ (.D(_01369_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[120][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15599_ (.D(_01370_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[120][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15600_ (.D(_01371_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[110][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15601_ (.D(_01372_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[110][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15602_ (.D(_01373_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[117][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15603_ (.D(_01374_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[117][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15604_ (.D(_01375_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[87][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15605_ (.D(_01376_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[87][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15606_ (.D(_01377_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[11][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15607_ (.D(_01378_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15608_ (.D(_01379_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[116][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15609_ (.D(_01380_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[116][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15610_ (.D(_01381_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[118][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15611_ (.D(_01382_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[118][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15612_ (.D(_01383_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[115][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15613_ (.D(_01384_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[115][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15614_ (.D(_01385_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[289][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15615_ (.D(_01386_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[289][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15616_ (.D(_01387_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[90][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15617_ (.D(_01388_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[90][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15618_ (.D(_01389_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[247][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15619_ (.D(_01390_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[247][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15620_ (.D(_01391_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15621_ (.D(_01392_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.bufreg2.i_cnt_done ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15622_ (.D(_01393_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.ctrl.i_jump ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15623_ (.D(_01394_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.mem_if.signbit ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15624_ (.D(_01395_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.state.genblk1.misalign_trap_sync_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15625_ (.D(_01396_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[88][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15626_ (.D(_01397_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[88][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15627_ (.D(_01398_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15628_ (.D(_01399_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15629_ (.D(_01400_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[279][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15630_ (.D(_01401_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[279][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15631_ (.D(_01402_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[244][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15632_ (.D(_01403_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[244][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15633_ (.D(_01404_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.state.o_cnt_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15634_ (.D(_01405_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.state.o_cnt_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15635_ (.D(_01406_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.state.o_cnt_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15636_ (.D(_01407_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.state.o_cnt_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15637_ (.D(_01408_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.state.o_cnt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15638_ (.D(_01409_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15639_ (.D(_01410_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15640_ (.D(_01411_),
    .CLK(net3),
    .Q(\mod.u_cpu.cpu.state.stage_two_req ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15641_ (.D(_01412_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[269][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15642_ (.D(_01413_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[269][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15643_ (.D(_01414_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[259][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15644_ (.D(_01415_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[259][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15645_ (.D(_01416_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[249][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _15646_ (.D(_01417_),
    .CLK(net3),
    .Q(\mod.u_cpu.rf_ram.memory[249][1] ));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_9 (.ZN(net9));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_10 (.ZN(net10));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_11 (.ZN(net11));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_12 (.ZN(net12));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_13 (.ZN(net13));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_14 (.ZN(net14));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_15 (.ZN(net15));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_16 (.ZN(net16));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_17 (.ZN(net17));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_18 (.ZN(net18));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_19 (.ZN(net19));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_20 (.ZN(net20));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_21 (.ZN(net21));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_22 (.ZN(net22));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_23 (.ZN(net23));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_24 (.ZN(net24));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_25 (.ZN(net25));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_26 (.ZN(net26));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_27 (.ZN(net27));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_28 (.ZN(net28));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_29 (.ZN(net29));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_30 (.ZN(net30));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_31 (.ZN(net31));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_32 (.ZN(net32));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_33 (.ZN(net33));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_34 (.ZN(net34));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_35 (.ZN(net35));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_36 (.ZN(net36));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_37 (.ZN(net37));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_38 (.ZN(net38));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_39 (.ZN(net39));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_40 (.ZN(net40));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_41 (.ZN(net41));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_42 (.ZN(net42));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_43 (.ZN(net43));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_44 (.ZN(net44));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_45 (.ZN(net45));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_46 (.ZN(net46));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_47 (.ZN(net47));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_48 (.ZN(net48));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_49 (.ZN(net49));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_50 (.ZN(net50));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_51 (.ZN(net51));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_52 (.ZN(net52));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_53 (.ZN(net53));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_54 (.ZN(net54));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_55 (.ZN(net55));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_56 (.ZN(net56));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_57 (.ZN(net57));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_58 (.ZN(net58));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_59 (.ZN(net59));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_60 (.ZN(net60));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_61 (.ZN(net61));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_62 (.ZN(net62));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_63 (.ZN(net63));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_64 (.ZN(net64));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_65 (.ZN(net65));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_66 (.ZN(net66));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_67 (.ZN(net67));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_68 (.ZN(net68));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_69 (.ZN(net69));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_70 (.ZN(net70));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_71 (.ZN(net71));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_72 (.ZN(net72));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_73 (.ZN(net73));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_74 (.ZN(net74));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_75 (.ZN(net75));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_76 (.ZN(net76));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_77 (.ZN(net77));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_78 (.ZN(net78));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_79 (.ZN(net79));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_80 (.ZN(net80));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_81 (.ZN(net81));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_82 (.ZN(net82));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_83 (.ZN(net83));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_84 (.ZN(net84));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_85 (.ZN(net85));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_86 (.ZN(net86));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_87 (.ZN(net87));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_88 (.ZN(net88));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_89 (.ZN(net89));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_90 (.ZN(net90));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_91 (.ZN(net91));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_92 (.ZN(net92));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_93 (.ZN(net93));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_94 (.ZN(net94));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_95 (.ZN(net95));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_96 (.ZN(net96));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_97 (.ZN(net97));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_98 (.ZN(net98));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_99 (.ZN(net99));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_100 (.ZN(net100));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_101 (.ZN(net101));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_102 (.ZN(net102));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_103 (.ZN(net103));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_104 (.ZN(net104));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_105 (.ZN(net105));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_106 (.ZN(net106));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_107 (.ZN(net107));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_108 (.ZN(net108));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_109 (.ZN(net109));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_110 (.ZN(net110));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_111 (.ZN(net111));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_112 (.ZN(net112));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_113 (.ZN(net113));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_114 (.ZN(net114));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_115 (.ZN(net115));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_116 (.ZN(net116));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_117 (.ZN(net117));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_118 (.ZN(net118));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_119 (.ZN(net119));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_120 (.ZN(net120));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_121 (.ZN(net121));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_122 (.ZN(net122));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_123 (.ZN(net123));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_124 (.ZN(net124));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_125 (.ZN(net125));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_126 (.ZN(net126));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_127 (.ZN(net127));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_128 (.ZN(net128));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_129 (.ZN(net129));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_130 (.ZN(net130));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_131 (.ZN(net131));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_132 (.ZN(net132));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_133 (.ZN(net133));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_134 (.ZN(net134));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_135 (.ZN(net135));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_136 (.ZN(net136));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_137 (.ZN(net137));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_138 (.ZN(net138));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_139 (.ZN(net139));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_140 (.ZN(net140));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_141 (.ZN(net141));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_142 (.ZN(net142));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_143 (.ZN(net143));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_144 (.ZN(net144));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_145 (.ZN(net145));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_146 (.ZN(net146));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_147 (.ZN(net147));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_148 (.ZN(net148));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_149 (.ZN(net149));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_150 (.ZN(net150));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_151 (.ZN(net151));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_152 (.ZN(net152));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_153 (.ZN(net153));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_154 (.ZN(net154));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_155 (.ZN(net155));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_156 (.ZN(net156));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_157 (.ZN(net157));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_158 (.ZN(net158));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_159 (.ZN(net159));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_160 (.ZN(net160));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_161 (.ZN(net161));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_162 (.ZN(net162));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_163 (.ZN(net163));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_164 (.ZN(net164));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_165 (.ZN(net165));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_166 (.ZN(net166));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_167 (.ZN(net167));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_168 (.ZN(net168));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_169 (.ZN(net169));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_170 (.ZN(net170));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_171 (.ZN(net171));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_172 (.ZN(net172));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_173 (.ZN(net173));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_174 (.ZN(net174));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_175 (.ZN(net175));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_176 (.ZN(net176));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_177 (.ZN(net177));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_178 (.ZN(net178));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_179 (.ZN(net179));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_180 (.ZN(net180));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_181 (.ZN(net181));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14224__D (.I(_00000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _15821_ (.I(net4),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_349 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_350 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_351 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_352 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_353 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_354 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_355 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_356 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_357 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_358 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_359 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_360 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_361 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_362 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_363 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_364 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_365 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_366 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_367 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_368 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_369 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_370 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_371 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_372 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_373 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_374 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_375 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_376 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_377 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_378 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_379 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_380 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_381 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_382 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_383 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_384 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_385 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_386 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_387 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_388 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_389 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_390 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_391 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_392 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_393 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_394 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_395 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_396 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_397 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_398 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_399 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_400 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_401 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_402 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_403 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_404 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_405 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_406 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_407 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_408 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_409 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_410 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_411 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_412 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_413 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_414 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_415 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_416 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_417 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_418 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_419 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_420 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_421 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_422 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_423 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_424 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_425 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_426 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_427 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_428 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_429 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_430 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_431 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_432 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_433 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_434 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_435 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_436 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_437 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_438 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_439 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_440 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_441 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_442 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_443 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_444 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_445 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_446 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_447 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_448 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_449 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_450 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_451 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_452 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_453 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_454 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_455 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_456 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_457 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_458 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_459 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_460 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_461 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_462 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_463 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_464 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_465 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_466 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_467 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_468 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_469 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_470 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_471 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_472 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_473 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_474 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_475 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_476 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_477 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_478 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_479 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_480 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_481 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_482 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_483 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_484 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_485 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_486 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_487 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_488 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_489 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_490 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_491 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_492 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_493 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_494 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_495 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_496 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_497 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_498 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_499 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_500 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_501 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_502 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_503 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_504 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_505 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_506 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_507 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_508 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_509 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_510 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_511 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_512 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_513 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_514 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_515 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_516 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_517 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_518 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_519 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_520 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_521 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_522 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_523 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_524 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_525 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_526 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_527 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_528 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_529 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_530 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_531 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_532 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5644 ();
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1 (.I(io_in[10]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(io_in[11]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__buf_20 input3 (.I(io_in[12]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 input4 (.I(io_in[8]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(io_in[9]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output6 (.I(net6),
    .Z(io_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output7 (.I(net7),
    .Z(io_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_8 (.ZN(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14225__D (.I(_00001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15312__D (.I(_00073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15240__D (.I(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15421__D (.I(_01196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15525__D (.I(_01296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15549__D (.I(_01320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15553__D (.I(_01324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09518__A1 (.I(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09491__S (.I(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09474__A1 (.I(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07110__A1 (.I(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08984__B (.I(_01421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08969__A1 (.I(_01421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08946__I (.I(_01421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07114__A1 (.I(_01421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08996__C (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08980__A4 (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08948__I (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07114__A2 (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12966__I (.I(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07146__C (.I(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07129__A1 (.I(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09025__A1 (.I(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09010__I (.I(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08981__A1 (.I(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07122__A1 (.I(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09009__A1 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09002__I (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08978__A1 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07122__A3 (.I(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09013__A1 (.I(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07143__A1 (.I(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07123__C (.I(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09477__A1 (.I(_01439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07151__I (.I(_01439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07139__I (.I(_01439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07132__A1 (.I(_01439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09479__B (.I(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08945__I (.I(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07142__A2 (.I(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07132__A2 (.I(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09498__I (.I(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09481__A2 (.I(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07134__B (.I(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07745__I (.I(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07732__I (.I(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07524__I (.I(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07136__I (.I(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08780__A1 (.I(_01446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07428__A1 (.I(_01446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07281__A1 (.I(_01446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07138__I (.I(_01446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08918__B (.I(_01447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08250__B (.I(_01447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08185__B (.I(_01447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07168__A1 (.I(_01447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09445__A1 (.I(_01451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07147__A2 (.I(_01451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09039__A2 (.I(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09031__A3 (.I(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07146__A1 (.I(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13899__A1 (.I(_01453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13004__A1 (.I(_01453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12979__A1 (.I(_01453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07145__A2 (.I(_01453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09494__A2 (.I(_01454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07146__A2 (.I(_01454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07540__I (.I(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07149__I (.I(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08938__A1 (.I(_01459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08415__A1 (.I(_01459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08275__A1 (.I(_01459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07168__A2 (.I(_01459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09523__B2 (.I(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09517__A1 (.I(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09480__A1 (.I(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07153__I (.I(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09507__A1 (.I(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09506__A1 (.I(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07164__A1 (.I(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07154__I (.I(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09951__A1 (.I(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07161__A1 (.I(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07159__A1 (.I(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07155__I (.I(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12857__A1 (.I(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08939__A1 (.I(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08276__A1 (.I(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07157__A1 (.I(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08939__A2 (.I(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08276__A2 (.I(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07158__A2 (.I(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07157__A2 (.I(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08860__A1 (.I(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07160__I (.I(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08606__A1 (.I(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07162__I (.I(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08859__A1 (.I(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08139__A1 (.I(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07729__A1 (.I(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07167__A2 (.I(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07430__I (.I(_01474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07166__I (.I(_01474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08858__A1 (.I(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08138__A1 (.I(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07839__B (.I(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07167__A3 (.I(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07169__I (.I(_01477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12845__A1 (.I(_01478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09832__A1 (.I(_01478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08943__S (.I(_01478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07173__A1 (.I(_01478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13756__A1 (.I(_01479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07173__A2 (.I(_01479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08744__B (.I(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08607__A1 (.I(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07973__B (.I(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07730__A1 (.I(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07840__I (.I(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07605__C (.I(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07175__I (.I(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08809__A1 (.I(_01483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08450__B (.I(_01483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08074__A1 (.I(_01483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07348__A1 (.I(_01483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07669__I (.I(_01484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07177__I (.I(_01484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08072__I (.I(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07731__I (.I(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07539__B (.I(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07178__I (.I(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08704__A1 (.I(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08626__A1 (.I(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07429__A1 (.I(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07282__A1 (.I(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07749__I (.I(_01487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07582__I (.I(_01487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07180__I (.I(_01487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08685__C (.I(_01489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08212__I (.I(_01489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07346__A1 (.I(_01489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07246__A1 (.I(_01489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07697__I (.I(_01491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07387__I (.I(_01491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07361__I (.I(_01491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07184__I (.I(_01491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08544__C (.I(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07294__I (.I(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07228__I (.I(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07185__I (.I(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08789__A1 (.I(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08037__A1 (.I(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07427__A1 (.I(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07227__A1 (.I(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09477__A2 (.I(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07336__I (.I(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07325__I (.I(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07187__I (.I(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08589__A1 (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08487__A1 (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08455__A1 (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07194__S0 (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07392__I (.I(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07260__I (.I(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07215__I (.I(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07190__I (.I(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07734__I (.I(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07546__I (.I(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07357__I (.I(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07192__I (.I(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08514__C (.I(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07247__S1 (.I(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07233__S1 (.I(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07194__S1 (.I(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07227__A2 (.I(_01502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07559__I (.I(_01503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07536__I (.I(_01503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07530__I (.I(_01503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07196__I (.I(_01503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08600__C (.I(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08543__C (.I(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07264__I (.I(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07197__I (.I(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07292__A1 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07257__A1 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07241__A1 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07222__A1 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08713__S0 (.I(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07632__A1 (.I(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07619__A1 (.I(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07200__I (.I(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08745__S (.I(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08291__S0 (.I(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07236__A1 (.I(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07206__A1 (.I(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07554__I (.I(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07402__I (.I(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07373__I (.I(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07202__I (.I(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07529__I (.I(_01510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07300__I (.I(_01510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07265__I (.I(_01510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07203__I (.I(_01510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08804__A1 (.I(_01511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07250__A1 (.I(_01511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07235__A1 (.I(_01511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07205__A1 (.I(_01511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10434__A1 (.I(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07205__A2 (.I(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07449__I (.I(_01515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07229__I (.I(_01515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07210__I (.I(_01515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07208__I (.I(_01515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08791__S (.I(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07892__A1 (.I(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07497__A1 (.I(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07218__A1 (.I(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08503__A1 (.I(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08483__A1 (.I(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07239__A1 (.I(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07214__A1 (.I(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10420__A1 (.I(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07214__A2 (.I(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08732__S1 (.I(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07256__C (.I(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07240__C (.I(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07218__C (.I(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07457__I (.I(_01527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07408__I (.I(_01527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07378__I (.I(_01527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07220__I (.I(_01527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08053__I (.I(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07343__I (.I(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07276__I (.I(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07221__I (.I(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07426__C (.I(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07257__C (.I(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07241__C (.I(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07222__C (.I(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08299__I (.I(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07983__I (.I(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07835__I (.I(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07226__I (.I(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08789__B (.I(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08037__B (.I(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07427__C (.I(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07227__C (.I(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08331__I (.I(_01537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07964__I (.I(_01537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07363__I (.I(_01537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07230__I (.I(_01537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08220__I (.I(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07396__I (.I(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07355__I (.I(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07231__I (.I(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07941__I (.I(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07299__I (.I(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07248__I (.I(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07232__I (.I(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08507__A1 (.I(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07285__S0 (.I(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07247__S0 (.I(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07233__S0 (.I(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08686__S (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07291__A1 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07256__A1 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07240__A1 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07562__I (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07411__I (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07369__I (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07243__I (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08069__I (.I(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07877__I (.I(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07310__I (.I(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07244__I (.I(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08839__S1 (.I(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08117__S1 (.I(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07258__C (.I(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07245__C (.I(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07258__A2 (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08694__I (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07435__I (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07270__I (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07253__I (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08798__S0 (.I(_01561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08363__A1 (.I(_01561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07290__A1 (.I(_01561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07255__A1 (.I(_01561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08668__A1 (.I(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08368__A1 (.I(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07399__A1 (.I(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07263__S0 (.I(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07818__I (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07438__I (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07329__I (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07261__I (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07998__I (.I(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07746__I (.I(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07463__I (.I(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07262__I (.I(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07313__S1 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07298__S1 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07285__S1 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07263__S1 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07280__A2 (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08700__A1 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07315__A1 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07287__A1 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07267__A1 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12528__A1 (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07267__A2 (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08840__S (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07319__A1 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07308__A1 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07275__A1 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08693__S0 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07318__A1 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07305__A1 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07272__A1 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08078__I (.I(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07702__I (.I(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07608__I (.I(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07274__I (.I(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07880__I (.I(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07319__C (.I(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07291__C (.I(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07275__C (.I(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08055__I (.I(_01586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07860__I (.I(_01586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07460__I (.I(_01586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07279__I (.I(_01586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08336__C (.I(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07321__C (.I(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07293__C (.I(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07280__C (.I(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08449__B (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08373__A1 (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08137__C (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07347__A1 (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08833__A1 (.I(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08346__A1 (.I(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08110__A1 (.I(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07312__A1 (.I(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07293__A2 (.I(_01593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08624__B (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07768__B (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07321__A1 (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07311__A1 (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07750__I (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07548__I (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07498__I (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07296__I (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07934__I (.I(_01604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07420__I (.I(_01604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07335__I (.I(_01604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07297__I (.I(_01604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08513__A1 (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07418__A1 (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07313__S0 (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07298__S0 (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07311__A2 (.I(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08293__A1 (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07911__A1 (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07334__A1 (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07303__A1 (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08853__A1 (.I(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08716__A1 (.I(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07333__A1 (.I(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07302__A1 (.I(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07308__B (.I(_01613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07959__I (.I(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07864__I (.I(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07424__I (.I(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07307__I (.I(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08452__I (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08334__C (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07342__C (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07308__C (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08797__B (.I(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08356__B (.I(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07345__C (.I(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07311__C (.I(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07321__A2 (.I(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08601__C (.I(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08468__C (.I(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07561__C (.I(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07324__I (.I(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08678__C (.I(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08615__B (.I(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07753__B (.I(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07345__A1 (.I(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07414__I (.I(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07389__I (.I(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07381__I (.I(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07326__I (.I(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08149__I (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07826__I (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07616__I (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07327__I (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08788__S0 (.I(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08278__I (.I(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08036__S0 (.I(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07331__S0 (.I(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08326__I (.I(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08042__I (.I(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07790__I (.I(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07330__I (.I(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08788__S1 (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08682__C (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08036__S1 (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07331__S1 (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07345__A2 (.I(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07640__A1 (.I(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07629__A1 (.I(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07615__A1 (.I(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07342__A1 (.I(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08098__I (.I(_01644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08061__I (.I(_01644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07655__I (.I(_01644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07337__I (.I(_01644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09474__A2 (.I(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07685__I (.I(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07444__I (.I(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07338__I (.I(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08102__I (.I(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07871__I (.I(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07853__I (.I(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07339__I (.I(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08847__S0 (.I(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08723__S0 (.I(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08711__S0 (.I(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07341__A1 (.I(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10149__A1 (.I(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07341__A2 (.I(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08344__C (.I(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08335__C (.I(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07916__A1 (.I(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07344__C (.I(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07509__A1 (.I(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08721__C (.I(_01657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07602__C (.I(_01657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07510__I (.I(_01657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07350__I (.I(_01657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08616__C (.I(_01658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08434__C (.I(_01658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08321__C (.I(_01658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07368__A1 (.I(_01658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09478__A1 (.I(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08457__I (.I(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07371__I (.I(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07353__I (.I(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07782__I (.I(_01661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07772__I (.I(_01661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07743__I (.I(_01661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07354__I (.I(_01661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08787__A1 (.I(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08611__B (.I(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08035__A1 (.I(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07360__A1 (.I(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08771__S0 (.I(_01664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08511__S (.I(_01664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08016__S0 (.I(_01664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07359__S0 (.I(_01664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08034__S1 (.I(_01666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07886__C (.I(_01666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07366__S1 (.I(_01666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07359__S1 (.I(_01666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07360__A2 (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08805__C (.I(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08701__C (.I(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07985__I (.I(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07362__I (.I(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08751__A1 (.I(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08646__A1 (.I(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07815__A1 (.I(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07367__A1 (.I(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07783__I (.I(_01671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07776__I (.I(_01671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07556__I (.I(_01671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07364__I (.I(_01671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08599__A1 (.I(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07817__I (.I(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07798__I (.I(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07365__I (.I(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08786__S0 (.I(_01673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08034__S0 (.I(_01673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07805__A1 (.I(_01673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07366__S0 (.I(_01673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07367__A2 (.I(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07769__I (.I(_01677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07593__C (.I(_01677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07528__I (.I(_01677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07370__I (.I(_01677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08425__C (.I(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08413__C (.I(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08312__C (.I(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07384__A1 (.I(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08353__I (.I(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08083__I (.I(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07525__I (.I(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07372__I (.I(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08749__C (.I(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08443__A1 (.I(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08437__A1 (.I(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07377__A1 (.I(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08773__A1 (.I(_01682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08201__I (.I(_01682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07885__A1 (.I(_01682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07376__S0 (.I(_01682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08533__C (.I(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07920__C (.I(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07382__S1 (.I(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07376__S1 (.I(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07377__A2 (.I(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07788__I (.I(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07664__I (.I(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07621__I (.I(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07379__I (.I(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08508__C (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08369__C (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07816__I (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07380__I (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08779__A1 (.I(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08234__I (.I(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08163__I (.I(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07383__A1 (.I(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07490__A1 (.I(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07476__A1 (.I(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07456__A1 (.I(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07382__S0 (.I(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07383__A2 (.I(_01690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07386__A2 (.I(_01692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08834__A1 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08111__A1 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08027__A1 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07386__B (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08854__C (.I(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08739__C (.I(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08730__C (.I(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07388__I (.I(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08785__A1 (.I(_01696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08665__C (.I(_01696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08033__A1 (.I(_01696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07413__A1 (.I(_01696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08574__A1 (.I(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08563__A1 (.I(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07663__A1 (.I(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07391__S0 (.I(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08720__A1 (.I(_01698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08590__C (.I(_01698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08456__C (.I(_01698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07391__S1 (.I(_01698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07413__A2 (.I(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07519__I (.I(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07474__I (.I(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07454__I (.I(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07393__I (.I(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07904__I (.I(_01701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07801__I (.I(_01701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07662__I (.I(_01701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07394__I (.I(_01701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08738__C (.I(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08729__C (.I(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08167__I (.I(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07395__I (.I(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08664__C (.I(_01703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08405__S1 (.I(_01703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07426__A1 (.I(_01703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07410__A1 (.I(_01703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08718__A1 (.I(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07758__I (.I(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07714__I (.I(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07397__I (.I(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08676__A1 (.I(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08186__I (.I(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07419__A1 (.I(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07400__A1 (.I(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08410__A1 (.I(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08400__A1 (.I(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08348__S (.I(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07407__A1 (.I(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07626__I (.I(_01710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07571__I (.I(_01710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07533__I (.I(_01710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07403__I (.I(_01710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08579__A1 (.I(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07705__A1 (.I(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07692__A1 (.I(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07405__A1 (.I(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08798__S1 (.I(_01714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08693__S1 (.I(_01714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07892__B (.I(_01714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07407__C (.I(_01714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08778__C (.I(_01717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08181__I (.I(_01717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08025__C (.I(_01717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07410__C (.I(_01717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08013__I (.I(_01719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07922__I (.I(_01719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07814__I (.I(_01719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07412__I (.I(_01719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08814__S1 (.I(_01720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08785__B (.I(_01720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08084__S1 (.I(_01720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07413__C (.I(_01720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08583__A1 (.I(_01722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07709__A1 (.I(_01722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07696__A1 (.I(_01722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07416__S0 (.I(_01722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08669__C (.I(_01723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08614__S1 (.I(_01723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07752__S1 (.I(_01723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07416__S1 (.I(_01723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07427__A2 (.I(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07487__A1 (.I(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07469__A1 (.I(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07448__A1 (.I(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07425__A1 (.I(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08494__A1 (.I(_01729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08474__A1 (.I(_01729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07716__A1 (.I(_01729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07423__A1 (.I(_01729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08847__S1 (.I(_01732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08723__S1 (.I(_01732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08711__S1 (.I(_01732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07425__C (.I(_01732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07426__B (.I(_01733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07428__A3 (.I(_01735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08658__B (.I(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08605__A1 (.I(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07728__A1 (.I(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07508__B (.I(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08857__C (.I(_01739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07971__A1 (.I(_01739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07668__A1 (.I(_01739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07507__A1 (.I(_01739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07948__A1 (.I(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07726__A1 (.I(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07667__A1 (.I(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07482__A1 (.I(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07862__I (.I(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07842__I (.I(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07462__I (.I(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07434__I (.I(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08320__C (.I(_01742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08311__C (.I(_01742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07969__A1 (.I(_01742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07461__A1 (.I(_01742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07733__I (.I(_01743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07611__I (.I(_01743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07517__I (.I(_01743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07436__I (.I(_01743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07990__I (.I(_01744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07822__I (.I(_01744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07466__I (.I(_01744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07437__I (.I(_01744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08176__I (.I(_01745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07600__A1 (.I(_01745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07484__S0 (.I(_01745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07440__S0 (.I(_01745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07910__I (.I(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07831__I (.I(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07763__I (.I(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07439__I (.I(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08229__I (.I(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08157__I (.I(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07484__S1 (.I(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07440__S1 (.I(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07461__A2 (.I(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07846__I (.I(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07652__I (.I(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07574__I (.I(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07442__I (.I(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07673__I (.I(_01750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07610__I (.I(_01750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07465__I (.I(_01750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07443__I (.I(_01750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08748__C (.I(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08319__C (.I(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08310__C (.I(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07459__A1 (.I(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07690__I (.I(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07654__I (.I(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07494__I (.I(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07445__I (.I(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08535__S0 (.I(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07493__S0 (.I(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07464__S0 (.I(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07447__A1 (.I(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08251__I (.I(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07718__I (.I(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07470__I (.I(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07450__I (.I(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07659__I (.I(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07641__I (.I(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07550__I (.I(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07451__I (.I(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07596__A1 (.I(_01759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07587__A1 (.I(_01759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07569__A1 (.I(_01759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07453__A1 (.I(_01759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08441__I (.I(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08359__I (.I(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07687__I (.I(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07455__I (.I(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08713__S1 (.I(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07534__S1 (.I(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07490__C (.I(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07456__C (.I(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08107__I (.I(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07858__I (.I(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07477__I (.I(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07458__I (.I(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07968__C (.I(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07956__C (.I(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07946__C (.I(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07459__C (.I(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07647__C (.I(_01768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07635__C (.I(_01768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07492__C (.I(_01768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07461__C (.I(_01768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08644__C (.I(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07811__C (.I(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07493__S1 (.I(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07464__S1 (.I(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07481__A2 (.I(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08422__C (.I(_01773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07503__A1 (.I(_01773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07491__A1 (.I(_01773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07478__A1 (.I(_01773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07637__S0 (.I(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07609__S0 (.I(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07486__A1 (.I(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07468__A1 (.I(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12533__A1 (.I(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07468__A2 (.I(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09517__A2 (.I(_01778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08103__I (.I(_01778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07872__I (.I(_01778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07471__I (.I(_01778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07894__I (.I(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07501__A1 (.I(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07489__A1 (.I(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07473__A1 (.I(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10567__A1 (.I(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07473__A2 (.I(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07633__C (.I(_01783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07620__C (.I(_01783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07502__C (.I(_01783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07476__C (.I(_01783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07775__I (.I(_01785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07503__C (.I(_01785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07491__C (.I(_01785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07478__C (.I(_01785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07899__I (.I(_01787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07699__I (.I(_01787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07504__I (.I(_01787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07480__I (.I(_01787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08593__B (.I(_01788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08517__B (.I(_01788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08460__B (.I(_01788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07481__C (.I(_01788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08566__A1 (.I(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07970__A1 (.I(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07636__A1 (.I(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07506__A1 (.I(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07492__A2 (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10531__A1 (.I(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07486__A2 (.I(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12429__A1 (.I(_01796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07489__A2 (.I(_01796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07505__A2 (.I(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08592__S0 (.I(_01802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08548__S0 (.I(_01802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07625__S0 (.I(_01802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07496__A1 (.I(_01802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07503__A2 (.I(_01805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08705__S (.I(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08679__S (.I(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08540__A1 (.I(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07502__A1 (.I(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10471__A1 (.I(_01808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07501__A2 (.I(_01808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08556__C (.I(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07666__C (.I(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07623__C (.I(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07505__C (.I(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07508__C (.I(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07730__A2 (.I(_01817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08631__A1 (.I(_01818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07781__A1 (.I(_01818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07754__C (.I(_01818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07527__A1 (.I(_01818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08132__A1 (.I(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07930__A1 (.I(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07855__A1 (.I(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07514__S0 (.I(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08051__I (.I(_01820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07856__I (.I(_01820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07522__I (.I(_01820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07513__I (.I(_01820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08343__C (.I(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07915__C (.I(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07516__S1 (.I(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07514__S1 (.I(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08091__A1 (.I(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08066__A1 (.I(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08050__A1 (.I(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07516__S0 (.I(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07630__I (.I(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07567__I (.I(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07535__I (.I(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07518__I (.I(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08537__S0 (.I(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07532__S0 (.I(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07523__S0 (.I(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07521__S0 (.I(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07944__I (.I(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07650__I (.I(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07624__I (.I(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07520__I (.I(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08133__C (.I(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08124__C (.I(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07532__S1 (.I(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07521__S1 (.I(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08830__C (.I(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08821__C (.I(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08106__C (.I(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07523__S1 (.I(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07526__I3 (.I(_01831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07670__I (.I(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07541__I (.I(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07538__S0 (.I(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07526__S0 (.I(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08534__C (.I(_01833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07887__C (.I(_01833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07538__S1 (.I(_01833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07526__S1 (.I(_01833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07527__A2 (.I(_01834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08878__C (.I(_01836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08636__A1 (.I(_01836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07793__A1 (.I(_01836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07539__A1 (.I(_01836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08594__S0 (.I(_01837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08461__S0 (.I(_01837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07545__S0 (.I(_01837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07531__S0 (.I(_01837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08461__S1 (.I(_01838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07584__S1 (.I(_01838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07545__S1 (.I(_01838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07531__S1 (.I(_01838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07538__I0 (.I(_01839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07538__I1 (.I(_01840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08518__S0 (.I(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08349__I (.I(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07594__S0 (.I(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07534__S0 (.I(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07538__I2 (.I(_01842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08539__A1 (.I(_01843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07584__S0 (.I(_01843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07565__S0 (.I(_01843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07537__S0 (.I(_01843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08518__S1 (.I(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07594__S1 (.I(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07565__S1 (.I(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07537__S1 (.I(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07538__I3 (.I(_01845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07539__A2 (.I(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08742__A1 (.I(_01848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08567__A1 (.I(_01848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08491__A1 (.I(_01848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07604__A1 (.I(_01848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08618__A1 (.I(_01849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08470__C (.I(_01849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07757__A1 (.I(_01849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07581__A1 (.I(_01849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09522__A1 (.I(_01850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07683__I (.I(_01850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07606__I (.I(_01850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07543__I (.I(_01850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08602__A1 (.I(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08469__A1 (.I(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07593__A1 (.I(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07563__A1 (.I(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07563__A2 (.I(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08786__S1 (.I(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08468__A1 (.I(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08235__I (.I(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07561__A1 (.I(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08784__S0 (.I(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08032__S0 (.I(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07723__A1 (.I(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07553__A1 (.I(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08596__A1 (.I(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08520__A1 (.I(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08463__A1 (.I(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07552__A1 (.I(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07995__I (.I(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07828__I (.I(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07808__I (.I(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07555__I (.I(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08776__A1 (.I(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08243__I (.I(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08023__A1 (.I(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07560__A1 (.I(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08523__A1 (.I(_01864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08466__A1 (.I(_01864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07986__I (.I(_01864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07558__A1 (.I(_01864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08524__C (.I(_01867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08467__C (.I(_01867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07591__C (.I(_01867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07560__C (.I(_01867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08740__C (.I(_01870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08712__B (.I(_01870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08500__C (.I(_01870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07563__C (.I(_01870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08670__C (.I(_01872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08526__A1 (.I(_01872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07602__A1 (.I(_01872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07580__A1 (.I(_01872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07580__A2 (.I(_01873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08525__A1 (.I(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07601__A1 (.I(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07592__A1 (.I(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07577__A1 (.I(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08498__A1 (.I(_01875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08478__A1 (.I(_01875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07597__A1 (.I(_01875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07570__A1 (.I(_01875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08524__A1 (.I(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08381__I (.I(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07591__A1 (.I(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07575__A1 (.I(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10913__A1 (.I(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07573__A2 (.I(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08290__I (.I(_01882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08044__I (.I(_01882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07600__C (.I(_01882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07575__C (.I(_01882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08545__I (.I(_01886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08370__I (.I(_01886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07681__I (.I(_01886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07579__I (.I(_01886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08602__C (.I(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08526__C (.I(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08469__C (.I(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07580__C (.I(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08856__C (.I(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08703__B (.I(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08547__B (.I(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07603__A1 (.I(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07593__A2 (.I(_01892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08612__S0 (.I(_01893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08521__A1 (.I(_01893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07747__S0 (.I(_01893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07588__A1 (.I(_01893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07602__A2 (.I(_01902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08423__I (.I(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07671__I (.I(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07648__I (.I(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07607__I (.I(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08777__C (.I(_01916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08535__S1 (.I(_01916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08024__C (.I(_01916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07609__S1 (.I(_01916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07623__A2 (.I(_01917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08432__C (.I(_01918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07646__A1 (.I(_01918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07634__A1 (.I(_01918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07622__A1 (.I(_01918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08444__I (.I(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08113__I (.I(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07649__I (.I(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07612__I (.I(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08501__S0 (.I(_01920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08492__S0 (.I(_01920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08481__S0 (.I(_01920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07614__A1 (.I(_01920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08623__S0 (.I(_01925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08171__I (.I(_01925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07767__S0 (.I(_01925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07620__A1 (.I(_01925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08592__S1 (.I(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08548__S1 (.I(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07637__S1 (.I(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07625__S1 (.I(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07635__A2 (.I(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08550__A1 (.I(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07675__A1 (.I(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07639__A1 (.I(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07628__A1 (.I(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08554__A1 (.I(_01938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07679__A1 (.I(_01938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07645__A1 (.I(_01938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07633__A1 (.I(_01938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08573__A1 (.I(_01949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08553__A1 (.I(_01949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07678__A1 (.I(_01949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07643__A1 (.I(_01949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08574__C (.I(_01952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08554__C (.I(_01952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07679__C (.I(_01952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07645__C (.I(_01952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08565__A1 (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08460__A1 (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07711__A1 (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07666__A1 (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08568__S0 (.I(_01957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08459__S0 (.I(_01957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07672__S0 (.I(_01957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07651__S0 (.I(_01957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08568__S1 (.I(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08459__S1 (.I(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07672__S1 (.I(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07651__S1 (.I(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07666__A2 (.I(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08564__A1 (.I(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08411__C (.I(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07710__A1 (.I(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07665__A1 (.I(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08570__A1 (.I(_01963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08559__A1 (.I(_01963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08360__S0 (.I(_01963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07657__A1 (.I(_01963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11387__A1 (.I(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07657__A2 (.I(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08604__A1 (.I(_01977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08528__A1 (.I(_01977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07924__A1 (.I(_01977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07727__A1 (.I(_01977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08741__A1 (.I(_01978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08586__A1 (.I(_01978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07923__C (.I(_01978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07701__A1 (.I(_01978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08593__A1 (.I(_01979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08576__A1 (.I(_01979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08402__C (.I(_01979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07682__A1 (.I(_01979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07682__A2 (.I(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08575__A1 (.I(_01981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08555__A1 (.I(_01981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08401__C (.I(_01981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07680__A1 (.I(_01981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11537__A1 (.I(_01982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07675__A2 (.I(_01982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14184__A1 (.I(_01985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07678__A2 (.I(_01985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08585__A1 (.I(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08412__C (.I(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07725__A1 (.I(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07700__A1 (.I(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08048__I (.I(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07896__I (.I(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07712__I (.I(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07686__I (.I(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08557__S0 (.I(_01994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08436__S0 (.I(_01994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07703__S0 (.I(_01994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07688__S0 (.I(_01994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08577__S1 (.I(_01995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08438__S1 (.I(_01995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07713__S1 (.I(_01995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07688__S1 (.I(_01995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07700__A2 (.I(_01996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08584__A1 (.I(_01997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08479__A1 (.I(_01997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07724__A1 (.I(_01997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07698__A1 (.I(_01997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08580__A1 (.I(_01998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08560__A1 (.I(_01998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07706__A1 (.I(_01998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07693__A1 (.I(_01998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08584__C (.I(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07724__C (.I(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07710__C (.I(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07698__C (.I(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08585__C (.I(_02007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08480__C (.I(_02007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07725__C (.I(_02007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07700__C (.I(_02007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08557__S1 (.I(_02010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08436__S1 (.I(_02010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08179__I (.I(_02010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07703__S1 (.I(_02010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07711__A2 (.I(_02011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11631__A1 (.I(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07705__A2 (.I(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08577__S0 (.I(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08442__S0 (.I(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08438__S0 (.I(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07713__S0 (.I(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07725__A2 (.I(_02021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08617__S0 (.I(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08475__A1 (.I(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07756__S0 (.I(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07717__A1 (.I(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07717__B (.I(_02024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08365__I (.I(_02026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07882__I (.I(_02026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07739__I (.I(_02026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07719__I (.I(_02026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08715__A1 (.I(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08582__A1 (.I(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08477__A1 (.I(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07721__A1 (.I(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08583__C (.I(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08478__C (.I(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08287__I (.I(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07723__C (.I(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07729__A3 (.I(_02036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07730__B (.I(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08899__A1 (.I(_02039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08323__A1 (.I(_02039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08214__A1 (.I(_02039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07771__A1 (.I(_02039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08609__A1 (.I(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08527__B (.I(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08302__I (.I(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07737__A1 (.I(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08504__A1 (.I(_02041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08495__A1 (.I(_02041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08484__A1 (.I(_02041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07736__S0 (.I(_02041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08739__A1 (.I(_02043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08730__A1 (.I(_02043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08617__S1 (.I(_02043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07736__S1 (.I(_02043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07737__A2 (.I(_02044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08620__A1 (.I(_02046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08603__B (.I(_02046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07761__A1 (.I(_02046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07744__A1 (.I(_02046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08627__S0 (.I(_02048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07881__S (.I(_02048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07773__S0 (.I(_02048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07742__S0 (.I(_02048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08610__S1 (.I(_02049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07898__C (.I(_02049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07773__S1 (.I(_02049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07742__S1 (.I(_02049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07744__A2 (.I(_02050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08783__A1 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08620__B (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07761__B (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07744__B (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08784__S1 (.I(_02054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08612__S1 (.I(_02054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08032__S1 (.I(_02054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07747__S1 (.I(_02054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08615__A1 (.I(_02057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08029__I (.I(_02057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07794__I (.I(_02057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07753__A1 (.I(_02057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08614__S0 (.I(_02059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08532__A1 (.I(_02059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08464__A1 (.I(_02059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07752__S0 (.I(_02059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07753__A2 (.I(_02060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08854__A1 (.I(_02063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08805__A1 (.I(_02063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08701__A1 (.I(_02063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07756__S1 (.I(_02063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08619__S0 (.I(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08296__A1 (.I(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07915__A1 (.I(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07760__S0 (.I(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08619__S1 (.I(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08608__S1 (.I(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08352__C (.I(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07760__S1 (.I(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07761__A2 (.I(_02068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08621__S0 (.I(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08597__A1 (.I(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07919__A1 (.I(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07764__S0 (.I(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08623__S1 (.I(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08621__S1 (.I(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07767__S1 (.I(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07764__S1 (.I(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07765__A2 (.I(_02072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08722__B (.I(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08624__A1 (.I(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08611__A1 (.I(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07768__A1 (.I(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07768__A2 (.I(_02075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08625__C (.I(_02077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08383__B (.I(_02077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08289__B (.I(_02077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07770__C (.I(_02077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07973__A1 (.I(_02079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12847__A1 (.I(_02080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08379__C (.I(_02080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08283__C (.I(_02080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07774__A1 (.I(_02080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07774__A2 (.I(_02081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08877__C (.I(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08393__A1 (.I(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08300__A1 (.I(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07780__A1 (.I(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08737__A1 (.I(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08728__A1 (.I(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08218__I (.I(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07777__I (.I(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08629__S0 (.I(_02085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08610__S0 (.I(_02085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08351__A1 (.I(_02085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07779__S0 (.I(_02085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08794__C (.I(_02086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08629__S1 (.I(_02086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08627__S1 (.I(_02086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07779__S1 (.I(_02086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08633__A1 (.I(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08628__A1 (.I(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08031__A1 (.I(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07787__A1 (.I(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08542__A1 (.I(_02091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07989__I (.I(_02091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07901__I (.I(_02091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07784__I (.I(_02091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08634__S0 (.I(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08632__S0 (.I(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07791__S0 (.I(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07786__S0 (.I(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08843__C (.I(_02093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08689__C (.I(_02093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08297__C (.I(_02093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07786__S1 (.I(_02093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08499__C (.I(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08488__C (.I(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08479__C (.I(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07789__I (.I(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08635__A1 (.I(_02097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08630__A1 (.I(_02097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08215__I (.I(_02097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07792__A1 (.I(_02097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08634__S1 (.I(_02098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08632__S1 (.I(_02098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08030__S1 (.I(_02098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07791__S1 (.I(_02098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08857__A1 (.I(_02102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08637__B (.I(_02102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08301__B (.I(_02102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07795__B (.I(_02102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07839__A1 (.I(_02103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08656__A1 (.I(_02105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08394__B (.I(_02105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08003__A1 (.I(_02105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07837__A1 (.I(_02105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08750__S0 (.I(_02106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08638__S0 (.I(_02106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08587__S (.I(_02106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07800__S0 (.I(_02106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08782__S1 (.I(_02107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08750__S1 (.I(_02107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08253__I (.I(_02107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07800__S1 (.I(_02107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07815__A2 (.I(_02108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08804__C (.I(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08368__C (.I(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08017__I (.I(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07802__I (.I(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08654__A1 (.I(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08645__A1 (.I(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07834__A1 (.I(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07813__A1 (.I(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08641__A1 (.I(_02111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08407__A1 (.I(_02111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08397__A1 (.I(_02111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07806__A1 (.I(_02111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07806__B (.I(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08644__A1 (.I(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08318__A1 (.I(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08153__I (.I(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07811__A1 (.I(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08643__A1 (.I(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08286__I (.I(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08154__I (.I(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07810__A1 (.I(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07813__B (.I(_02119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08231__I (.I(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08159__I (.I(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07921__A1 (.I(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07813__C (.I(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08655__A1 (.I(_02124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08141__I (.I(_02124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07984__A1 (.I(_02124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07836__A1 (.I(_02124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08647__S0 (.I(_02125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08453__S (.I(_02125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07974__S0 (.I(_02125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07820__S0 (.I(_02125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08085__I (.I(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08080__I (.I(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07844__I (.I(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07819__I (.I(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08647__S1 (.I(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08638__S1 (.I(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07974__S1 (.I(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07820__S1 (.I(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07836__A2 (.I(_02128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08650__A1 (.I(_02129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08148__I (.I(_02129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07978__A1 (.I(_02129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07825__A1 (.I(_02129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07825__B (.I(_02132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08653__A1 (.I(_02135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08047__A1 (.I(_02135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07981__A1 (.I(_02135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07832__A1 (.I(_02135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08652__A1 (.I(_02136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08600__A1 (.I(_02136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07980__A1 (.I(_02136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07830__A1 (.I(_02136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08653__C (.I(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08270__I (.I(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07981__C (.I(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07832__C (.I(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08654__C (.I(_02141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08645__C (.I(_02141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07982__C (.I(_02141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07834__C (.I(_02141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08655__C (.I(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08440__A1 (.I(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08161__I (.I(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07836__C (.I(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07837__A3 (.I(_02144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07838__A2 (.I(_02145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08743__C (.I(_02148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08529__A1 (.I(_02148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08374__A1 (.I(_02148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07972__A1 (.I(_02148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08761__B (.I(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08136__A1 (.I(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08071__A1 (.I(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07879__A1 (.I(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08832__A1 (.I(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08135__A1 (.I(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08109__A1 (.I(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07861__A1 (.I(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08835__S0 (.I(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08127__S0 (.I(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07925__S0 (.I(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07845__S0 (.I(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08835__S1 (.I(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08143__I (.I(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08112__S1 (.I(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07845__S1 (.I(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07861__A2 (.I(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08719__C (.I(_02154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08097__I (.I(_02154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07866__I (.I(_02154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07847__I (.I(_02154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08384__S1 (.I(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08134__A1 (.I(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07932__A1 (.I(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07859__A1 (.I(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08747__A1 (.I(_02156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08242__I (.I(_02156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08130__A1 (.I(_02156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07852__A1 (.I(_02156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08129__A1 (.I(_02157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07927__A1 (.I(_02157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07869__A1 (.I(_02157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07851__A1 (.I(_02157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08793__A1 (.I(_02161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08726__A1 (.I(_02161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08133__A1 (.I(_02161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07857__A1 (.I(_02161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12750__A1 (.I(_02162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07855__A2 (.I(_02162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08537__S1 (.I(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07931__C (.I(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07875__C (.I(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07857__C (.I(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08134__C (.I(_02166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07932__C (.I(_02166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07876__C (.I(_02166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07859__C (.I(_02166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08126__C (.I(_02168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07957__C (.I(_02168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07933__C (.I(_02168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07861__C (.I(_02168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08813__S0 (.I(_02171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08754__A1 (.I(_02171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08082__S0 (.I(_02171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07865__S0 (.I(_02171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07949__S1 (.I(_02172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07935__S1 (.I(_02172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07925__S1 (.I(_02172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07865__S1 (.I(_02172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07878__A2 (.I(_02173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07968__A1 (.I(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07956__A1 (.I(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07946__A1 (.I(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07876__A1 (.I(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08175__I (.I(_02175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07952__A1 (.I(_02175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07928__A1 (.I(_02175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07870__A1 (.I(_02175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08735__A1 (.I(_02179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08688__A1 (.I(_02179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07931__A1 (.I(_02179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07875__A1 (.I(_02179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07966__A1 (.I(_02180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07954__A1 (.I(_02180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07943__A1 (.I(_02180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07874__A1 (.I(_02180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12149__A1 (.I(_02181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07874__A2 (.I(_02181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08823__C (.I(_02185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08135__C (.I(_02185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08094__C (.I(_02185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07878__C (.I(_02185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07924__A2 (.I(_02187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08534__A1 (.I(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08392__A1 (.I(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08282__C (.I(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07887__A1 (.I(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07887__A2 (.I(_02189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08852__A1 (.I(_02190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08803__A1 (.I(_02190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08699__A1 (.I(_02190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07883__I (.I(_02190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08843__A1 (.I(_02191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08391__A1 (.I(_02191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08297__A1 (.I(_02191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07886__A1 (.I(_02191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11928__A1 (.I(_02192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07886__A2 (.I(_02192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07886__B (.I(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08546__A1 (.I(_02196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08392__C (.I(_02196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08298__C (.I(_02196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07900__A1 (.I(_02196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08734__A1 (.I(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08725__A1 (.I(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08333__A1 (.I(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07890__I (.I(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08319__A1 (.I(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08310__A1 (.I(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08281__A1 (.I(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07893__A1 (.I(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12745__A1 (.I(_02199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07893__A2 (.I(_02199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08794__A1 (.I(_02202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08689__A1 (.I(_02202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08673__A1 (.I(_02202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07898__A1 (.I(_02202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11970__A1 (.I(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07898__A2 (.I(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08801__A1 (.I(_02204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08758__A1 (.I(_02204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08697__A1 (.I(_02204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07897__A1 (.I(_02204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07898__B (.I(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07900__A3 (.I(_02206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08536__B (.I(_02207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07969__C (.I(_02207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07947__C (.I(_02207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07900__B (.I(_02207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08708__A1 (.I(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08199__I (.I(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08142__I (.I(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07906__A1 (.I(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08811__S0 (.I(_02211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08796__S0 (.I(_02211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08752__S0 (.I(_02211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07905__A1 (.I(_02211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08853__C (.I(_02212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08700__C (.I(_02212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07975__I (.I(_02212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07905__B (.I(_02212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08543__A1 (.I(_02216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08226__I (.I(_02216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08192__I (.I(_02216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07909__A1 (.I(_02216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08837__S1 (.I(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08347__I (.I(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08115__S1 (.I(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07911__C (.I(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08757__A1 (.I(_02220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08385__I (.I(_02220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08342__A1 (.I(_02220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07914__A1 (.I(_02220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11999__A1 (.I(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07914__A2 (.I(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08533__A1 (.I(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08416__S0 (.I(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08315__A1 (.I(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07920__A1 (.I(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12046__A1 (.I(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07920__A2 (.I(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07923__B1 (.I(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08751__B (.I(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08684__A1 (.I(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08447__A1 (.I(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07923__B2 (.I(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07933__A2 (.I(_02233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12808__A1 (.I(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07927__A2 (.I(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08838__S0 (.I(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08116__S0 (.I(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07949__S0 (.I(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07935__S0 (.I(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07947__A2 (.I(_02243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08431__A1 (.I(_02244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08421__A1 (.I(_02244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07963__A1 (.I(_02244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07940__A1 (.I(_02244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08258__I (.I(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07962__A1 (.I(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07951__A1 (.I(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07939__A1 (.I(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08782__S0 (.I(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08030__S0 (.I(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07955__A1 (.I(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07945__A1 (.I(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08594__S1 (.I(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07967__C (.I(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07955__C (.I(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07945__C (.I(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07957__A2 (.I(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08812__S0 (.I(_02266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08081__S0 (.I(_02266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08046__A1 (.I(_02266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07960__S0 (.I(_02266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08813__S1 (.I(_02267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08116__S1 (.I(_02267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08082__S1 (.I(_02267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07960__S1 (.I(_02267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07969__A2 (.I(_02268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08842__A1 (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08530__S (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08390__A1 (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07967__A1 (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07972__A3 (.I(_02279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07973__C (.I(_02280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07984__A2 (.I(_02282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08769__A1 (.I(_02283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08012__A1 (.I(_02283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08001__A1 (.I(_02283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07982__A1 (.I(_02283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13107__A1 (.I(_02284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07977__A2 (.I(_02284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07982__B (.I(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08779__C (.I(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08210__I (.I(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08026__C (.I(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07984__C (.I(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08770__A1 (.I(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08026__A1 (.I(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08014__A1 (.I(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08002__A1 (.I(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08762__S0 (.I(_02294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08666__S (.I(_02294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08004__S0 (.I(_02294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07988__S0 (.I(_02294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08762__S1 (.I(_02295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08544__A1 (.I(_02295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08004__S1 (.I(_02295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07988__S1 (.I(_02295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08002__A2 (.I(_02296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08765__A1 (.I(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08020__A1 (.I(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08007__A1 (.I(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07993__A1 (.I(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08764__A1 (.I(_02298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08019__A1 (.I(_02298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08006__A1 (.I(_02298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07992__A1 (.I(_02298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08818__A1 (.I(_02302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08089__A1 (.I(_02302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08064__A1 (.I(_02302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07999__A1 (.I(_02302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08767__A1 (.I(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08467__A1 (.I(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08010__A1 (.I(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07997__A1 (.I(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08768__C (.I(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08207__I (.I(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08011__C (.I(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07999__C (.I(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08769__C (.I(_02308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08247__I (.I(_02308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08012__C (.I(_02308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08001__C (.I(_02308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08028__A2 (.I(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08014__A2 (.I(_02312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08827__A1 (.I(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08768__A1 (.I(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08101__A1 (.I(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08011__A1 (.I(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08770__C (.I(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08183__I (.I(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08033__B (.I(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08014__C (.I(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08027__A2 (.I(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08771__S1 (.I(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08601__A1 (.I(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08391__C (.I(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08016__S1 (.I(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08778__A1 (.I(_02325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08416__S1 (.I(_02325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08237__I (.I(_02325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08025__A1 (.I(_02325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08777__A1 (.I(_02329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08164__I (.I(_02329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08121__A1 (.I(_02329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08024__A1 (.I(_02329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12224__A1 (.I(_02330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08023__A2 (.I(_02330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08025__B (.I(_02332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08026__B (.I(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08808__A1 (.I(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08449__A1 (.I(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08137__A1 (.I(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08073__A1 (.I(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08038__A1 (.I(_02339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08035__A2 (.I(_02342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08038__B2 (.I(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08073__A2 (.I(_02346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08720__C (.I(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08324__I (.I(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08057__I (.I(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08040__I (.I(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08797__A1 (.I(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08692__A1 (.I(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08094__A1 (.I(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08056__A1 (.I(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08845__S0 (.I(_02349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08691__S0 (.I(_02349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08086__S0 (.I(_02349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08043__S0 (.I(_02349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08691__S1 (.I(_02350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08304__I (.I(_02350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08114__S1 (.I(_02350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08043__S1 (.I(_02350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08056__A2 (.I(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08759__A1 (.I(_02352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08093__A1 (.I(_02352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08068__A1 (.I(_02352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08054__A1 (.I(_02352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13061__A1 (.I(_02353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08046__A2 (.I(_02353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08054__A2 (.I(_02355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08850__A1 (.I(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08092__A1 (.I(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08067__A1 (.I(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08052__A1 (.I(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08758__C (.I(_02359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08092__C (.I(_02359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08067__C (.I(_02359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08052__C (.I(_02359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08759__C (.I(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08093__C (.I(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08068__C (.I(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08054__C (.I(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08832__C (.I(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08760__C (.I(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08109__C (.I(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08056__C (.I(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08846__A1 (.I(_02365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08823__A1 (.I(_02365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08126__A1 (.I(_02365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08070__A1 (.I(_02365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08815__S0 (.I(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08810__S0 (.I(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08076__S0 (.I(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08060__S0 (.I(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08824__S1 (.I(_02367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08815__S1 (.I(_02367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08096__S1 (.I(_02367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08060__S1 (.I(_02367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08070__A2 (.I(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08817__A1 (.I(_02369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08115__S0 (.I(_02369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08088__A1 (.I(_02369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08063__A1 (.I(_02369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13049__A1 (.I(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08066__A2 (.I(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08068__B (.I(_02375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08846__B (.I(_02377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08692__B (.I(_02377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08345__C (.I(_02377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08070__C (.I(_02377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08073__B (.I(_02379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08834__C (.I(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08808__C (.I(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08111__C (.I(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08073__C (.I(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08810__S1 (.I(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08127__S1 (.I(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08118__S1 (.I(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08076__S1 (.I(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08707__A1 (.I(_02385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08355__S0 (.I(_02385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08337__S0 (.I(_02385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08079__S0 (.I(_02385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08811__S1 (.I(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08796__S1 (.I(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08752__S1 (.I(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08079__S1 (.I(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08838__S1 (.I(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08812__S1 (.I(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08165__I (.I(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08081__S1 (.I(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08084__I2 (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08084__I3 (.I(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08839__S0 (.I(_02391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08814__S0 (.I(_02391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08117__S0 (.I(_02391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08084__S0 (.I(_02391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08111__A2 (.I(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08845__S1 (.I(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08836__S1 (.I(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08187__I (.I(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08086__S1 (.I(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08094__A2 (.I(_02394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08089__B (.I(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08824__S0 (.I(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08118__S0 (.I(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08112__S0 (.I(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08096__S0 (.I(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08109__A2 (.I(_02404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08831__A1 (.I(_02405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08822__A1 (.I(_02405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08125__A1 (.I(_02405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08108__A1 (.I(_02405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08837__S0 (.I(_02406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08826__A1 (.I(_02406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08120__A1 (.I(_02406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08100__A1 (.I(_02406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08108__A2 (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08830__A1 (.I(_02410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08821__A1 (.I(_02410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08124__A1 (.I(_02410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08106__A1 (.I(_02410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08829__A1 (.I(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08820__A1 (.I(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08123__A1 (.I(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08105__A1 (.I(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11746__A1 (.I(_02412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08105__A2 (.I(_02412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08831__C (.I(_02415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08822__C (.I(_02415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08125__C (.I(_02415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08108__C (.I(_02415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08138__A2 (.I(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08117__I0 (.I(_02420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08836__S0 (.I(_02421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08339__A1 (.I(_02421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08329__A1 (.I(_02421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08114__S0 (.I(_02421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08117__I1 (.I(_02422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08117__I2 (.I(_02423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08117__I3 (.I(_02424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08137__A2 (.I(_02425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08126__A2 (.I(_02426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08135__A2 (.I(_02435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10398__A1 (.I(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08129__A2 (.I(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08134__A2 (.I(_02438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10263__A1 (.I(_02439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08132__A2 (.I(_02439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08137__B (.I(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08908__A1 (.I(_02449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08888__A1 (.I(_02449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08198__A1 (.I(_02449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08162__A1 (.I(_02449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08861__S0 (.I(_02450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08661__A1 (.I(_02450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08264__S0 (.I(_02450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08144__S0 (.I(_02450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08880__S1 (.I(_02451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08861__S1 (.I(_02451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08264__S1 (.I(_02451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08144__S1 (.I(_02451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08162__A2 (.I(_02452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08507__C (.I(_02453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08498__C (.I(_02453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08487__C (.I(_02453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08146__I (.I(_02453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08313__S1 (.I(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08303__S1 (.I(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08217__I (.I(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08147__I (.I(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08887__A1 (.I(_02455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08868__A1 (.I(_02455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08196__A1 (.I(_02455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08160__A1 (.I(_02455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08883__A1 (.I(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08864__A1 (.I(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08191__A1 (.I(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08152__A1 (.I(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08889__S0 (.I(_02457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08882__A1 (.I(_02457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08190__A1 (.I(_02457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08151__A1 (.I(_02457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08886__A1 (.I(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08867__A1 (.I(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08195__A1 (.I(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08158__A1 (.I(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08866__A1 (.I(_02462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08677__A1 (.I(_02462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08408__A1 (.I(_02462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08156__A1 (.I(_02462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08886__C (.I(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08795__A1 (.I(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08195__C (.I(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08158__C (.I(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08907__C (.I(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08887__C (.I(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08196__C (.I(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08160__C (.I(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08908__C (.I(_02469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08263__C (.I(_02469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08233__C (.I(_02469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08162__C (.I(_02469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08917__A1 (.I(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08897__A1 (.I(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08211__A1 (.I(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08184__A1 (.I(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08870__S0 (.I(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08863__A1 (.I(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08266__A1 (.I(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08166__S0 (.I(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08889__S1 (.I(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08870__S1 (.I(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08200__S1 (.I(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08166__S1 (.I(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08184__A2 (.I(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08426__S1 (.I(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08395__S1 (.I(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08382__S1 (.I(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08168__I (.I(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08774__A1 (.I(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08682__A1 (.I(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08238__I (.I(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08170__I (.I(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08891__A1 (.I(_02479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08872__A1 (.I(_02479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08674__A1 (.I(_02479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08173__A1 (.I(_02479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08895__C (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08876__C (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08298__A1 (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08180__C (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08916__C (.I(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08896__C (.I(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08209__C (.I(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08182__C (.I(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08917__C (.I(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08273__C (.I(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08249__C (.I(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08184__C (.I(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08185__A2 (.I(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08900__S0 (.I(_02494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08880__S0 (.I(_02494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08216__S0 (.I(_02494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08188__S0 (.I(_02494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08919__S1 (.I(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08900__S1 (.I(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08216__S1 (.I(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08188__S1 (.I(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08198__A2 (.I(_02496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08196__A2 (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08905__A1 (.I(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08885__A1 (.I(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08398__A1 (.I(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08194__A1 (.I(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12850__A1 (.I(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08927__C (.I(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08888__C (.I(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08198__C (.I(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08909__S0 (.I(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08902__A1 (.I(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08236__S0 (.I(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08200__S0 (.I(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08211__A2 (.I(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08930__A1 (.I(_02509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08911__A1 (.I(_02509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08240__A1 (.I(_02509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08203__A1 (.I(_02509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08934__C (.I(_02515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08915__C (.I(_02515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08246__C (.I(_02515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08208__C (.I(_02515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08936__C (.I(_02518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08897__C (.I(_02518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08869__C (.I(_02518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08211__C (.I(_02518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08937__B (.I(_02520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08898__B (.I(_02520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08274__B (.I(_02520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08213__B (.I(_02520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08276__A3 (.I(_02522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12849__A1 (.I(_02523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08927__A1 (.I(_02523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08263__A1 (.I(_02523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08233__A1 (.I(_02523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08233__A2 (.I(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08514__A1 (.I(_02526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08428__A1 (.I(_02526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08418__A1 (.I(_02526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08219__I (.I(_02526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08922__A1 (.I(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08903__A1 (.I(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08257__A1 (.I(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08223__A1 (.I(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08928__S0 (.I(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08921__A1 (.I(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08256__A1 (.I(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08222__A1 (.I(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08755__A1 (.I(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08387__A1 (.I(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08309__A1 (.I(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08225__I (.I(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08924__A1 (.I(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08429__A1 (.I(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08419__A1 (.I(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08228__A1 (.I(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08926__C (.I(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08413__A1 (.I(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08262__C (.I(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08232__C (.I(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08936__A1 (.I(_02542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08869__A1 (.I(_02542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08273__A1 (.I(_02542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08249__A1 (.I(_02542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08928__S1 (.I(_02543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08909__S1 (.I(_02543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08678__A1 (.I(_02543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08236__S1 (.I(_02543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08249__A2 (.I(_02544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08931__A1 (.I(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08912__A1 (.I(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08267__A1 (.I(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08241__A1 (.I(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08934__A1 (.I(_02550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08915__A1 (.I(_02550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08271__A1 (.I(_02550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08246__A1 (.I(_02550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08933__A1 (.I(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08914__A1 (.I(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08269__A1 (.I(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08245__A1 (.I(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09941__A1 (.I(_02552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08245__A2 (.I(_02552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08935__C (.I(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08868__C (.I(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08272__C (.I(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08248__C (.I(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08384__S0 (.I(_02559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08340__A1 (.I(_02559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08330__A1 (.I(_02559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08252__I (.I(_02559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08919__S0 (.I(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08378__A1 (.I(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08282__A1 (.I(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08254__S0 (.I(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08665__A1 (.I(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08379__A1 (.I(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08283__A1 (.I(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08254__S1 (.I(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08263__A2 (.I(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08664__A1 (.I(_02566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08316__A1 (.I(_02566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08307__A1 (.I(_02566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08260__A1 (.I(_02566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08273__A2 (.I(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08867__C (.I(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08844__A1 (.I(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08690__A1 (.I(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08271__C (.I(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08277__B (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08748__A1 (.I(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08375__S (.I(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08294__A1 (.I(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08279__S (.I(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08283__A2 (.I(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08721__A1 (.I(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08683__C (.I(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08380__I (.I(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08285__I (.I(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08878__A1 (.I(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08321__A1 (.I(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08312__A1 (.I(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08289__A1 (.I(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08313__S0 (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08306__A1 (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08303__S0 (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08288__S0 (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08709__A1 (.I(_02594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08683__A1 (.I(_02594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08378__C (.I(_02594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08288__S1 (.I(_02594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08289__A2 (.I(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08677__C (.I(_02597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08344__A1 (.I(_02597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08335__A1 (.I(_02597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08291__S1 (.I(_02597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08300__A2 (.I(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08297__B (.I(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08671__A1 (.I(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08403__C (.I(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08393__C (.I(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08300__C (.I(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08879__B (.I(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08435__A1 (.I(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08414__A1 (.I(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08322__A1 (.I(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08312__A2 (.I(_02610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08749__A1 (.I(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08424__A1 (.I(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08320__A1 (.I(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08311__A1 (.I(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08311__A2 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08321__A2 (.I(_02620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08316__B (.I(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08318__A2 (.I(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08760__A1 (.I(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08356__A1 (.I(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08345__A1 (.I(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08336__A1 (.I(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08738__A1 (.I(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08729__A1 (.I(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08681__A1 (.I(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08327__S0 (.I(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08708__C (.I(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08355__S1 (.I(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08337__S1 (.I(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08327__S1 (.I(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08336__A2 (.I(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08335__A2 (.I(_02637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08608__S0 (.I(_02638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08364__A1 (.I(_02638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08343__A1 (.I(_02638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08334__A1 (.I(_02638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08333__A2 (.I(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08345__A2 (.I(_02644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08342__A2 (.I(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08345__B (.I(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08433__A1 (.I(_02654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08412__A1 (.I(_02654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08402__A1 (.I(_02654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08354__A1 (.I(_02654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08354__A2 (.I(_02655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08660__A1 (.I(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08411__A1 (.I(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08377__A1 (.I(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08352__A1 (.I(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08352__B (.I(_02658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08844__C (.I(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08795__C (.I(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08690__C (.I(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08354__C (.I(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08356__A2 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08807__C (.I(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08510__A1 (.I(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08490__A1 (.I(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08372__B (.I(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08806__A1 (.I(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08702__A1 (.I(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08509__A1 (.I(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08371__A1 (.I(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08501__S1 (.I(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08492__S1 (.I(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08481__S1 (.I(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08360__S1 (.I(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08371__A2 (.I(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08508__A1 (.I(_02668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08499__A1 (.I(_02668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08488__A1 (.I(_02668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08369__A1 (.I(_02668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08369__A2 (.I(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08506__A1 (.I(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08497__A1 (.I(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08486__A1 (.I(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08367__A1 (.I(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08367__A2 (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08806__C (.I(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08509__C (.I(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08489__C (.I(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08371__C (.I(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08372__C (.I(_02678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08379__A2 (.I(_02682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08590__A1 (.I(_02688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08426__S0 (.I(_02688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08395__S0 (.I(_02688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08382__S0 (.I(_02688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08383__A2 (.I(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08393__A2 (.I(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08391__B (.I(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08403__A2 (.I(_02702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08397__A2 (.I(_02703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08403__B (.I(_02709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08669__A1 (.I(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08663__A1 (.I(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08456__A1 (.I(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08405__S0 (.I(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08413__A2 (.I(_02712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08407__A2 (.I(_02713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08536__A1 (.I(_02730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08446__A1 (.I(_02730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08433__C (.I(_02730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08424__C (.I(_02730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08434__A2 (.I(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08428__A2 (.I(_02734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08450__A1 (.I(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08437__A2 (.I(_02743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08439__A2 (.I(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08516__S1 (.I(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08472__S1 (.I(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08445__S1 (.I(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08442__S1 (.I(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08443__A2 (.I(_02749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08719__A1 (.I(_02751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08516__S0 (.I(_02751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08472__S0 (.I(_02751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08445__S0 (.I(_02751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08446__A2 (.I(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08449__A2 (.I(_02755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08450__A2 (.I(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08607__A2 (.I(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08670__A1 (.I(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08591__A1 (.I(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08515__A1 (.I(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08458__A1 (.I(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08458__A2 (.I(_02760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08458__B (.I(_02763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08709__C (.I(_02764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08591__C (.I(_02764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08515__C (.I(_02764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08458__C (.I(_02764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08460__A2 (.I(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08469__A2 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08491__A2 (.I(_02777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08480__A2 (.I(_02779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08479__A2 (.I(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08477__A2 (.I(_02783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08489__A2 (.I(_02788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08500__A2 (.I(_02799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08497__A2 (.I(_02803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08509__A2 (.I(_02808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08506__A2 (.I(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08515__A2 (.I(_02818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08515__B (.I(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08517__A2 (.I(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08526__A2 (.I(_02825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08520__A2 (.I(_02826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08525__A2 (.I(_02828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08523__A2 (.I(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08534__A2 (.I(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08536__A2 (.I(_02842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08546__A2 (.I(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08542__A2 (.I(_02848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08855__C (.I(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08731__C (.I(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08702__C (.I(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08546__C (.I(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08556__A2 (.I(_02855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08565__A2 (.I(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08567__A3 (.I(_02873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08576__A2 (.I(_02875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08570__A2 (.I(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08573__A2 (.I(_02879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08585__A2 (.I(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08604__A2 (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08591__A2 (.I(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08593__A2 (.I(_02899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08602__A2 (.I(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08601__A2 (.I(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08599__A2 (.I(_02905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08607__B (.I(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08609__A2 (.I(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08611__A2 (.I(_02917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08615__A2 (.I(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08620__A2 (.I(_02926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08622__A2 (.I(_02928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08624__A2 (.I(_02930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08744__A1 (.I(_02933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08628__A2 (.I(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08630__A2 (.I(_02936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08658__A1 (.I(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08645__B (.I(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08655__A2 (.I(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08650__B (.I(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08656__A3 (.I(_02962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08657__A2 (.I(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08660__A2 (.I(_02966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08663__A2 (.I(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08669__A2 (.I(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08678__A2 (.I(_02981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08676__A2 (.I(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08683__A2 (.I(_02986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08682__B (.I(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08743__A1 (.I(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08690__A2 (.I(_02993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08689__B (.I(_02995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08692__A2 (.I(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08703__A2 (.I(_02999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08702__A2 (.I(_03000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08849__A1 (.I(_03001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08800__A1 (.I(_03001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08732__S0 (.I(_03001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08696__A1 (.I(_03001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08701__A2 (.I(_03004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08699__A2 (.I(_03005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08704__A2 (.I(_03010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08709__A2 (.I(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08708__A2 (.I(_03013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08709__B (.I(_03015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08855__A1 (.I(_03017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08740__A1 (.I(_03017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08731__A1 (.I(_03017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08712__A1 (.I(_03017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08712__A2 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08722__A2 (.I(_03019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08721__A2 (.I(_03020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08720__A2 (.I(_03023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08718__A2 (.I(_03024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08731__A2 (.I(_03030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08740__A2 (.I(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08734__A2 (.I(_03040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08737__A2 (.I(_03043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08742__A3 (.I(_03048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08761__A1 (.I(_03056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08751__A2 (.I(_03057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08760__A2 (.I(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08770__A2 (.I(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08780__A2 (.I(_03077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08776__A2 (.I(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08778__B (.I(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08779__B (.I(_03085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08809__A2 (.I(_03088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08783__A2 (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08787__A2 (.I(_03093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08808__A2 (.I(_03097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08794__B (.I(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08797__A2 (.I(_03103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08806__A2 (.I(_03105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08805__A2 (.I(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08803__A2 (.I(_03109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08808__B (.I(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08814__I1 (.I(_03118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08814__I2 (.I(_03119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08814__I3 (.I(_03120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08834__A2 (.I(_03121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08823__A2 (.I(_03122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08817__A2 (.I(_03123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08822__A2 (.I(_03125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08832__A2 (.I(_03131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08831__A2 (.I(_03134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08829__A2 (.I(_03135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08858__A2 (.I(_03141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08839__I0 (.I(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08839__I1 (.I(_03143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08839__I2 (.I(_03144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08839__I3 (.I(_03145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08857__A2 (.I(_03146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08844__A2 (.I(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08856__A1 (.I(_03151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08846__A2 (.I(_03152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08855__A2 (.I(_03154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08856__B (.I(_03162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08869__A2 (.I(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08878__A2 (.I(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08878__B (.I(_03184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08888__A2 (.I(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08887__A2 (.I(_03190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08897__A2 (.I(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08899__A3 (.I(_03205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08908__A2 (.I(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08917__A2 (.I(_03216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08927__A2 (.I(_03226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08921__A2 (.I(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08936__A2 (.I(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08940__B (.I(_03246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13506__A2 (.I(_03250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09050__I (.I(_03250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09048__A1 (.I(_03250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09047__C (.I(_03250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09028__B (.I(_03251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08992__I (.I(_03251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08976__A1 (.I(_03251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08947__I (.I(_03251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08988__B (.I(_03256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08973__A1 (.I(_03256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08952__I (.I(_03256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09040__A3 (.I(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09036__A2 (.I(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09018__A1 (.I(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08955__A2 (.I(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13509__A3 (.I(_03260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09009__A3 (.I(_03260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08991__A1 (.I(_03260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09450__A3 (.I(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08961__A2 (.I(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13932__A1 (.I(_03268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12978__I (.I(_03268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09023__B (.I(_03268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08972__A1 (.I(_03268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13932__C (.I(_03269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12977__I (.I(_03269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09023__A2 (.I(_03269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08965__A1 (.I(_03269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14159__A2 (.I(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08972__A2 (.I(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13317__A1 (.I(_03271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09523__A1 (.I(_03271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08967__A2 (.I(_03271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09463__A2 (.I(_03276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08998__I0 (.I(_03276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08972__B (.I(_03276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13932__B (.I(_03279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09117__I (.I(_03279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09092__B2 (.I(_03279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08988__A1 (.I(_03279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12453__A1 (.I(_03289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09437__A1 (.I(_03289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08986__A1 (.I(_03289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13532__I (.I(_03292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09465__I (.I(_03292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09011__A2 (.I(_03292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08988__A2 (.I(_03292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13641__A1 (.I(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13640__A1 (.I(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09093__I (.I(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09014__A1 (.I(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14164__A1 (.I(_03298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13762__A1 (.I(_03298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09021__A1 (.I(_03298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09014__A2 (.I(_03298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09092__B1 (.I(_03300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09065__A1 (.I(_03300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08996__B (.I(_03300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13509__A2 (.I(_03302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09029__I (.I(_03302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08998__I1 (.I(_03302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13611__B (.I(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09013__A2 (.I(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13901__A1 (.I(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09058__A1 (.I(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09023__A1 (.I(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09006__A1 (.I(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14068__I (.I(_03309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13607__A1 (.I(_03309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09007__A2 (.I(_03309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09005__A2 (.I(_03309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13508__A2 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09043__A1 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09025__B (.I(_03329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13838__A1 (.I(_03331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09440__A2 (.I(_03331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09439__I (.I(_03331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09028__C (.I(_03331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13838__B (.I(_03334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09448__A1 (.I(_03334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09075__I (.I(_03334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09032__A1 (.I(_03334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12986__A2 (.I(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09032__A2 (.I(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13514__B (.I(_03337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12991__B1 (.I(_03337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09460__A2 (.I(_03337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09037__A1 (.I(_03337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12967__A1 (.I(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12861__I (.I(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12459__A1 (.I(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09035__A1 (.I(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12980__A2 (.I(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09040__A4 (.I(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09042__B (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09455__A1 (.I(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09094__I (.I(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09047__A1 (.I(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09046__A1 (.I(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09507__A2 (.I(_03352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09049__I (.I(_03352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13001__A2 (.I(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12973__B2 (.I(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09444__A1 (.I(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09067__A1 (.I(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13903__A1 (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12461__A2 (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09064__B1 (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09057__A1 (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13902__A1 (.I(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12461__A1 (.I(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12459__B (.I(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09057__C (.I(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13605__A1 (.I(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09123__A1 (.I(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09092__A1 (.I(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09064__A1 (.I(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14162__A1 (.I(_03363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09133__A1 (.I(_03363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09122__A1 (.I(_03363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09064__A2 (.I(_03363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13714__A1 (.I(_03364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13699__A1 (.I(_03364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09064__B2 (.I(_03364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09066__A2 (.I(_03368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12970__I (.I(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09067__A2 (.I(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13428__A1 (.I(_03371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09446__A1 (.I(_03371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09227__A1 (.I(_03371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09073__A1 (.I(_03371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09592__A1 (.I(_03374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09495__A1 (.I(_03374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09489__A2 (.I(_03374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09072__I (.I(_03374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13770__B (.I(_03377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13422__A1 (.I(_03377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12465__A3 (.I(_03377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09076__I (.I(_03377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13614__A2 (.I(_03378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13613__A1 (.I(_03378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09081__A2 (.I(_03378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09080__A1 (.I(_03378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09102__A1 (.I(_03383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09123__A2 (.I(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09109__I (.I(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09100__A1 (.I(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09085__I (.I(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09397__A1 (.I(_03386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09368__A1 (.I(_03386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09341__A1 (.I(_03386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09086__I (.I(_03386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09138__A2 (.I(_03387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09134__A2 (.I(_03387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09131__A2 (.I(_03387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09102__A2 (.I(_03387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14199__A1 (.I(_03389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14194__A2 (.I(_03389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12975__A1 (.I(_03389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09089__A3 (.I(_03389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13933__B (.I(_03390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13643__A1 (.I(_03390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13258__A1 (.I(_03390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09090__I (.I(_03390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13767__A2 (.I(_03391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13383__A2 (.I(_03391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09443__I (.I(_03391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09096__A2 (.I(_03391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09129__I (.I(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09124__A1 (.I(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09119__A2 (.I(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09092__A2 (.I(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09102__B1 (.I(_03397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12852__I (.I(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09106__A1 (.I(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09098__A1 (.I(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09397__B1 (.I(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09368__B1 (.I(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09341__B1 (.I(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09101__I (.I(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09430__A2 (.I(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09347__B1 (.I(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09324__B1 (.I(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09102__B2 (.I(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13919__A1 (.I(_03403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13770__A1 (.I(_03403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09441__A2 (.I(_03403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09104__I (.I(_03403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13838__A2 (.I(_03404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12997__A2 (.I(_03404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09112__A1 (.I(_03404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12462__A2 (.I(_03406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09223__I (.I(_03406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09107__A2 (.I(_03406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09304__I (.I(_03407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09258__I (.I(_03407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09108__I (.I(_03407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09353__B1 (.I(_03408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09253__B1 (.I(_03408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09244__C1 (.I(_03408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09112__A2 (.I(_03408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09229__A1 (.I(_03410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09220__A1 (.I(_03410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09137__A2 (.I(_03410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09111__A1 (.I(_03410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13970__A1 (.I(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13170__A2 (.I(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12447__A1 (.I(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09120__A1 (.I(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09313__I (.I(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09164__I (.I(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09118__I (.I(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09115__I (.I(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09236__A1 (.I(_03414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09212__I (.I(_03414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09203__I (.I(_03414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09116__I (.I(_03414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09353__A1 (.I(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09317__A1 (.I(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09125__A2 (.I(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09120__A2 (.I(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09429__A1 (.I(_03417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09382__B (.I(_03417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09150__I (.I(_03417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09119__B (.I(_03417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13735__A2 (.I(_03424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13280__A2 (.I(_03424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12951__A2 (.I(_03424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09131__A1 (.I(_03424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13749__A2 (.I(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13289__A2 (.I(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09134__A1 (.I(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09347__A1 (.I(_03436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09324__A1 (.I(_03436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09157__A2 (.I(_03436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09143__A2 (.I(_03436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13956__B2 (.I(_03438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13952__B (.I(_03438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13949__A1 (.I(_03438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09147__I1 (.I(_03438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09419__A1 (.I(_03439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09412__A1 (.I(_03439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09405__A1 (.I(_03439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09147__S (.I(_03439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09162__S (.I(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09159__S (.I(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09154__S (.I(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09151__S (.I(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13968__B2 (.I(_03444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13963__A1 (.I(_03444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13960__A1 (.I(_03444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09154__I1 (.I(_03444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13991__A1 (.I(_03449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13789__I1 (.I(_03449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13389__A2 (.I(_03449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09162__I0 (.I(_03449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09194__I (.I(_03451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09185__I (.I(_03451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09176__I (.I(_03451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09165__I (.I(_03451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14007__A1 (.I(_03456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13229__I1 (.I(_03456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13191__A2 (.I(_03456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09173__I0 (.I(_03456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14012__A1 (.I(_03458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13633__I1 (.I(_03458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12943__A2 (.I(_03458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09177__I0 (.I(_03458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09183__S (.I(_03459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09181__S (.I(_03459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09179__S (.I(_03459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09177__S (.I(_03459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09201__S (.I(_03469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09199__S (.I(_03469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09197__S (.I(_03469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09195__S (.I(_03469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09210__S (.I(_03474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09208__S (.I(_03474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09206__S (.I(_03474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09204__S (.I(_03474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09253__A1 (.I(_03479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09217__S (.I(_03479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09215__S (.I(_03479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09213__S (.I(_03479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09228__A1 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09352__B (.I(_03488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09294__I (.I(_03488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09272__I (.I(_03488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09226__I (.I(_03488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09373__A1 (.I(_03489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09363__A1 (.I(_03489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09359__A1 (.I(_03489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09227__A2 (.I(_03489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09430__B1 (.I(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09396__B (.I(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09246__I (.I(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09232__A2 (.I(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09303__I (.I(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09280__I (.I(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09257__I (.I(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09235__I (.I(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09421__A1 (.I(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09392__A1 (.I(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09374__A1 (.I(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09244__A1 (.I(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09319__I (.I(_03497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09244__B1 (.I(_03497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12945__I (.I(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12443__I (.I(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09263__A4 (.I(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09238__I (.I(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13183__A1 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12947__A1 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12942__A1 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09240__I (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13789__S (.I(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13227__I (.I(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09249__I (.I(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09242__I (.I(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13872__A1 (.I(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13633__S (.I(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09255__A3 (.I(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09243__A2 (.I(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09271__A1 (.I(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09266__A1 (.I(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09261__A1 (.I(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09254__A1 (.I(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13816__S (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13750__A1 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13171__A1 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09251__A2 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09372__B1 (.I(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09362__B1 (.I(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09281__I (.I(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09259__I (.I(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09284__A3 (.I(_03521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09268__A2 (.I(_03521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09264__A2 (.I(_03521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09293__A1 (.I(_03528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09287__A1 (.I(_03528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09283__A1 (.I(_03528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09276__A1 (.I(_03528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09299__A1 (.I(_03535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09292__A1 (.I(_03535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09286__A1 (.I(_03535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09282__A1 (.I(_03535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09299__B1 (.I(_03536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09292__B1 (.I(_03536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09286__B1 (.I(_03536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09282__B1 (.I(_03536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09345__A2 (.I(_03538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09322__A2 (.I(_03538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09290__A2 (.I(_03538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09285__A2 (.I(_03538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09358__A1 (.I(_03554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09334__A1 (.I(_03554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09329__A1 (.I(_03554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09305__A1 (.I(_03554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09358__B1 (.I(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09334__B1 (.I(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09329__B1 (.I(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09305__B1 (.I(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09425__A2 (.I(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09411__A2 (.I(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09409__A1 (.I(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09312__C (.I(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09317__B1 (.I(_03562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09385__I (.I(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09372__A1 (.I(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09362__A1 (.I(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09316__A1 (.I(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09423__A1 (.I(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09390__A1 (.I(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09382__A1 (.I(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09315__A2 (.I(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09369__A1 (.I(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09348__A1 (.I(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09342__A1 (.I(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09325__A1 (.I(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09379__A3 (.I(_03586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09356__A2 (.I(_03586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09342__A3 (.I(_03586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09351__A1 (.I(_03590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09349__A2 (.I(_03590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09346__A2 (.I(_03590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13970__A2 (.I(_03614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09417__A1 (.I(_03614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09403__A1 (.I(_03614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09376__I (.I(_03614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09418__A2 (.I(_03615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09404__A2 (.I(_03615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09391__A2 (.I(_03615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09383__A2 (.I(_03615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13490__A1 (.I(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13486__B2 (.I(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09380__A1 (.I(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09378__B (.I(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09382__A2 (.I(_03617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13496__A1 (.I(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13494__B2 (.I(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09416__A3 (.I(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09400__A1 (.I(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09424__A4 (.I(_03637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09402__I (.I(_03637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13599__B2 (.I(_03659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13597__A1 (.I(_03659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09430__A1 (.I(_03659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13384__A1 (.I(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13365__I1 (.I(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10973__A1 (.I(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09442__A1 (.I(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13365__I0 (.I(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13322__A1 (.I(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09490__A1 (.I(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09435__A3 (.I(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13383__A1 (.I(_03665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11666__A1 (.I(_03665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10034__A2 (.I(_03665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09435__A4 (.I(_03665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13422__A2 (.I(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12459__A2 (.I(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09448__A2 (.I(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09438__I (.I(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13598__A2 (.I(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13520__A2 (.I(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12933__A2 (.I(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09442__B (.I(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14165__A1 (.I(_03670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13832__A2 (.I(_03670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13769__A1 (.I(_03670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09441__A1 (.I(_03670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13383__A3 (.I(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13258__A2 (.I(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09442__C (.I(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14194__B1 (.I(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13768__A1 (.I(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09445__A2 (.I(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09444__B (.I(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13425__A2 (.I(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12867__A1 (.I(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09451__B (.I(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09449__B (.I(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13910__A1 (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13832__B (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09461__A2 (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09453__A2 (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13908__A1 (.I(_03681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13640__A2 (.I(_03681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09461__A1 (.I(_03681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09455__A2 (.I(_03681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13835__A2 (.I(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13834__C (.I(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09457__A3 (.I(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09456__A4 (.I(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13761__A1 (.I(_03686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12995__I (.I(_03686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12464__C (.I(_03686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09462__A1 (.I(_03686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13611__A2 (.I(_03687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09462__A2 (.I(_03687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13587__I (.I(_03692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13578__I (.I(_03692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13569__I (.I(_03692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09466__I (.I(_03692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13599__A1 (.I(_03694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13597__A2 (.I(_03694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13596__A2 (.I(_03694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09468__B (.I(_03694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09551__I (.I(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09513__I (.I(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09470__I (.I(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12314__I (.I(_03696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11749__I (.I(_03696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09741__I (.I(_03696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09471__I (.I(_03696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09901__I (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09766__I (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09708__I (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09472__I (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12720__I (.I(_03698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12208__I (.I(_03698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11931__I (.I(_03698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09473__I (.I(_03698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14218__I0 (.I(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14213__I0 (.I(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14188__I0 (.I(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09504__I1 (.I(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12451__A1 (.I(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09569__A1 (.I(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09558__A1 (.I(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09475__A2 (.I(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09546__I (.I(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09476__I (.I(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09996__A1 (.I(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09704__A1 (.I(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09629__A1 (.I(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09486__A1 (.I(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09609__A1 (.I(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09484__A1 (.I(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09751__A1 (.I(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09733__A1 (.I(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09723__A1 (.I(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09486__A2 (.I(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12158__I (.I(_03712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11408__I (.I(_03712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09487__I (.I(_03712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13600__A1 (.I(_03713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13075__A1 (.I(_03713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10601__I (.I(_03713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09488__I (.I(_03713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10407__A1 (.I(_03714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09975__A1 (.I(_03714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09744__A1 (.I(_03714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09503__A1 (.I(_03714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10035__A2 (.I(_03715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09529__I (.I(_03715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09523__A2 (.I(_03715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09490__A2 (.I(_03715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10035__A3 (.I(_03717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09530__A2 (.I(_03717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09492__A2 (.I(_03717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09593__A1 (.I(_03718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09496__A1 (.I(_03718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10380__A1 (.I(_03721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10268__A1 (.I(_03721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09531__A2 (.I(_03721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09496__A2 (.I(_03721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10120__A1 (.I(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09951__A2 (.I(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09497__I (.I(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12691__A1 (.I(_03723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11604__A1 (.I(_03723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10774__A1 (.I(_03723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09502__A1 (.I(_03723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10973__A3 (.I(_03724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10859__A3 (.I(_03724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09703__A1 (.I(_03724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09499__A3 (.I(_03724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09594__A1 (.I(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09500__I (.I(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12234__A1 (.I(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12159__A1 (.I(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10395__A1 (.I(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09502__A2 (.I(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12702__A1 (.I(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12034__A1 (.I(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09503__A2 (.I(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09511__S (.I(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09504__S (.I(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11450__I (.I(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09538__I (.I(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09508__I (.I(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11632__I (.I(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10606__I (.I(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09747__I (.I(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09509__I (.I(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13078__I (.I(_03734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12773__I (.I(_03734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12688__I (.I(_03734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09510__I (.I(_03734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14220__I0 (.I(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14215__I0 (.I(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09712__I1 (.I(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09511__I1 (.I(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11235__I (.I(_03737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10740__I (.I(_03737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10193__I (.I(_03737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09514__I (.I(_03737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10053__I (.I(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09912__I (.I(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09731__I (.I(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09515__I (.I(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09683__I (.I(_03739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09645__I (.I(_03739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09588__I (.I(_03739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09516__I (.I(_03739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09583__I0 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09575__I0 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09564__I0 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09536__I0 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09760__A1 (.I(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09568__A2 (.I(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09525__A2 (.I(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11918__I (.I(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11076__I (.I(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09527__I (.I(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13235__A1 (.I(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12819__A1 (.I(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10267__I (.I(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09528__I (.I(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11335__A2 (.I(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10048__A1 (.I(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09844__A1 (.I(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09535__A1 (.I(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11839__A3 (.I(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10162__A2 (.I(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10034__A3 (.I(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09532__A1 (.I(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09831__A1 (.I(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09531__A1 (.I(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12272__A1 (.I(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11276__A1 (.I(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10465__A1 (.I(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09532__A2 (.I(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09544__I (.I(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09533__I (.I(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09815__A1 (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09655__I (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09602__I (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09534__I (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09582__A1 (.I(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09574__A1 (.I(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09563__A1 (.I(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09535__A2 (.I(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10996__I (.I(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10555__I (.I(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10095__I (.I(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09539__I (.I(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09971__I (.I(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09864__I (.I(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09698__I (.I(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09540__I (.I(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09577__I0 (.I(_03764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09566__I0 (.I(_03764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09556__I0 (.I(_03764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09542__I0 (.I(_03764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09772__I (.I(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09714__I (.I(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09628__I (.I(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09545__I (.I(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11992__A1 (.I(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09823__A1 (.I(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09614__A1 (.I(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09550__A1 (.I(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11284__I (.I(_03769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10277__I (.I(_03769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09548__I (.I(_03769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12825__A1 (.I(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12391__A1 (.I(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12049__I (.I(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09549__I (.I(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13241__A1 (.I(_03771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12063__A2 (.I(_03771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09849__A1 (.I(_03771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09550__A2 (.I(_03771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12005__I (.I(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11486__I (.I(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10619__I (.I(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09552__I (.I(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14208__A1 (.I(_03775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09633__A1 (.I(_03775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09615__A1 (.I(_03775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09554__A1 (.I(_03775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11939__I (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11087__I (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09561__I (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13246__A1 (.I(_03781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12830__A1 (.I(_03781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10287__I (.I(_03781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09562__I (.I(_03781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11457__A2 (.I(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10060__A1 (.I(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09854__A1 (.I(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09563__A2 (.I(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09874__A2 (.I(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09589__A2 (.I(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09579__A2 (.I(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09571__A1 (.I(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09797__A1 (.I(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09723__A2 (.I(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09647__A1 (.I(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09571__A2 (.I(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13407__A1 (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12743__A1 (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10495__I (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09573__I (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11522__A2 (.I(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10293__A1 (.I(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10065__A1 (.I(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09574__A2 (.I(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11952__I (.I(_03795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11100__I (.I(_03795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09580__I (.I(_03795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14144__A1 (.I(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12602__A1 (.I(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10298__I (.I(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09581__I (.I(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11582__A2 (.I(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10071__A1 (.I(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09868__A1 (.I(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09582__A2 (.I(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09617__I0 (.I(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09606__I0 (.I(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09600__I0 (.I(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09586__I0 (.I(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09641__I0 (.I(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09623__I0 (.I(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09604__I0 (.I(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09598__I0 (.I(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11711__I (.I(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10904__I (.I(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09590__I (.I(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14171__A1 (.I(_03804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14095__A1 (.I(_03804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10084__I (.I(_03804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09591__I (.I(_03804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11648__A2 (.I(_03805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09882__A1 (.I(_03805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09603__A2 (.I(_03805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09597__A1 (.I(_03805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09830__I (.I(_03806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09593__A2 (.I(_03806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10395__A2 (.I(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09702__I (.I(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09594__A2 (.I(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11144__A1 (.I(_03809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09859__I (.I(_03809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09684__I (.I(_03809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09596__I (.I(_03809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09606__S (.I(_03815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09604__S (.I(_03815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09936__A1 (.I(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09828__A2 (.I(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09762__A1 (.I(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09611__A1 (.I(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11321__I (.I(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10090__I (.I(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09612__I (.I(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14182__A1 (.I(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14149__A1 (.I(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09685__I (.I(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09613__I (.I(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14110__A1 (.I(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11744__A2 (.I(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09888__A1 (.I(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09614__A2 (.I(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12016__I (.I(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10917__I (.I(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09620__I (.I(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14127__A1 (.I(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13007__A1 (.I(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10100__I (.I(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09621__I (.I(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11821__A2 (.I(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09895__A1 (.I(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09781__A2 (.I(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09622__A2 (.I(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09653__I0 (.I(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09643__I0 (.I(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09635__I0 (.I(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09626__I0 (.I(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12004__A1 (.I(_03834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11987__A1 (.I(_03834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09765__A1 (.I(_03834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09632__A1 (.I(_03834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14105__A1 (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14088__A1 (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09860__I (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09631__I (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13012__A1 (.I(_03837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11945__A2 (.I(_03837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09900__A1 (.I(_03837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09632__A2 (.I(_03837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12079__I (.I(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10929__I (.I(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09638__I (.I(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14187__A1 (.I(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14122__A1 (.I(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10113__I (.I(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09639__I (.I(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12122__A2 (.I(_03843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09925__A2 (.I(_03843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09907__A1 (.I(_03843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09640__A2 (.I(_03843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12368__I (.I(_03849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11347__I (.I(_03849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09648__I (.I(_03849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14132__A1 (.I(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12105__A1 (.I(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10342__I (.I(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09649__I (.I(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12029__A2 (.I(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09986__A2 (.I(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09914__A1 (.I(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09650__A2 (.I(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11725__I (.I(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10942__I (.I(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09658__I (.I(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14072__A1 (.I(_03858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13054__A1 (.I(_03858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10129__I (.I(_03858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09659__I (.I(_03858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12285__A2 (.I(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10055__A2 (.I(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09920__A1 (.I(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09660__A2 (.I(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09664__S (.I(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09661__S (.I(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14083__A1 (.I(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12737__A1 (.I(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10354__I (.I(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09668__I (.I(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12374__A2 (.I(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11810__A2 (.I(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10136__A1 (.I(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09669__A2 (.I(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09672__S (.I(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09670__S (.I(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09820__A1 (.I(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09787__A1 (.I(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09715__A1 (.I(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09675__A1 (.I(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11736__I (.I(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10954__I (.I(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09676__I (.I(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13892__A1 (.I(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12754__A1 (.I(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10141__I (.I(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09677__I (.I(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12503__A2 (.I(_03873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10198__A2 (.I(_03873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09931__A1 (.I(_03873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09678__A2 (.I(_03873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09681__S (.I(_03874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09679__S (.I(_03874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09727__I0 (.I(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09719__I0 (.I(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09696__I0 (.I(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09687__I0 (.I(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13093__A2 (.I(_03878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12058__A2 (.I(_03878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09781__A1 (.I(_03878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09686__A1 (.I(_03878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12620__A1 (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12333__A1 (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11122__A1 (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09686__A2 (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09689__S (.I(_03880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09687__S (.I(_03880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11752__I (.I(_03884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10967__I (.I(_03884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09693__I (.I(_03884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14100__A1 (.I(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12726__A1 (.I(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10154__I (.I(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09694__I (.I(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12631__A2 (.I(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10328__A2 (.I(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09946__A1 (.I(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09695__A2 (.I(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09838__I (.I(_03889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09793__I (.I(_03889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09757__I (.I(_03889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09699__I (.I(_03889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09739__I0 (.I(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09729__I0 (.I(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09721__I0 (.I(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09700__I0 (.I(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11932__A1 (.I(_03892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11384__A1 (.I(_03892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10602__A1 (.I(_03892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09703__A2 (.I(_03892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11974__A1 (.I(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09744__A2 (.I(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09707__A1 (.I(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14207__A1 (.I(_03895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12684__A1 (.I(_03895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10773__I (.I(_03895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09706__I (.I(_03895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10396__A2 (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10167__A1 (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09952__A1 (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09707__A2 (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09712__S (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09711__A2 (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09710__A2 (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11027__I (.I(_03898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10432__I (.I(_03898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10168__I (.I(_03898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09709__I (.I(_03898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13601__I1 (.I(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10000__A1 (.I(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09953__A1 (.I(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09710__A1 (.I(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09754__A1 (.I(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09736__A1 (.I(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09726__A1 (.I(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09718__A1 (.I(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11771__I (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10980__I (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09716__I (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13030__A1 (.I(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12697__A1 (.I(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10173__I (.I(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09717__I (.I(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12796__A2 (.I(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10453__A2 (.I(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09957__A1 (.I(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09718__A2 (.I(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12184__I (.I(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11192__I (.I(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09724__I (.I(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14077__A1 (.I(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13412__A1 (.I(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10180__I (.I(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09725__I (.I(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14117__A2 (.I(_03911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10519__A2 (.I(_03911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09962__A1 (.I(_03911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09726__A2 (.I(_03911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09873__I (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09841__I (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09786__I (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09732__I (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09782__I0 (.I(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09777__I0 (.I(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09755__I0 (.I(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09737__I0 (.I(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11784__I (.I(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10992__I (.I(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09734__I (.I(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13064__A1 (.I(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12715__A1 (.I(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10186__I (.I(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09735__I (.I(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13018__A2 (.I(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10578__A2 (.I(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09968__A1 (.I(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09736__A2 (.I(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11228__I (.I(_03924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10796__I (.I(_03924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10406__I (.I(_03924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09743__I (.I(_03924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10025__I1 (.I(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09976__I1 (.I(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09816__I1 (.I(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09745__I1 (.I(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09749__S (.I(_03926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09745__S (.I(_03926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14174__I (.I(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10386__I (.I(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10002__I (.I(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09748__I (.I(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09978__I1 (.I(_03929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09955__I1 (.I(_03929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09818__I1 (.I(_03929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09749__I1 (.I(_03929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11797__I (.I(_03931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11008__I (.I(_03931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09752__I (.I(_03931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13082__A1 (.I(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12732__A1 (.I(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10203__I (.I(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09753__I (.I(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14177__A2 (.I(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10701__A2 (.I(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09981__A1 (.I(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09754__A2 (.I(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09784__I0 (.I(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09779__I0 (.I(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09770__I0 (.I(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09758__I0 (.I(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13120__A1 (.I(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13087__A1 (.I(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10810__I (.I(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09764__I (.I(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11826__A2 (.I(_03942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10418__A1 (.I(_03942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10209__A1 (.I(_03942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09765__A2 (.I(_03942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09770__S (.I(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09769__A2 (.I(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09768__A2 (.I(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12685__I (.I(_03944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12236__I (.I(_03944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11766__I (.I(_03944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09767__I (.I(_03944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09889__A1 (.I(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09850__A1 (.I(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09836__A1 (.I(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09768__A1 (.I(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11815__I (.I(_03949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11020__I (.I(_03949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09774__I (.I(_03949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13098__A1 (.I(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12765__A1 (.I(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10214__I (.I(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09775__I (.I(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11853__A2 (.I(_03951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10822__A2 (.I(_03951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09991__A1 (.I(_03951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09776__A2 (.I(_03951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11833__I (.I(_03959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11033__I (.I(_03959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09788__I (.I(_03959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13110__A1 (.I(_03960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12776__A1 (.I(_03960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10228__I (.I(_03960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09789__I (.I(_03960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10949__A2 (.I(_03961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10123__A2 (.I(_03961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10005__A1 (.I(_03961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09790__A2 (.I(_03961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09820__A2 (.I(_03966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09813__A2 (.I(_03966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09805__A2 (.I(_03966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09797__A2 (.I(_03966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12247__I (.I(_03967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11243__I (.I(_03967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09798__I (.I(_03967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14212__A1 (.I(_03968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12881__A1 (.I(_03968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10235__I (.I(_03968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09799__I (.I(_03968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11015__A2 (.I(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10760__A2 (.I(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10013__A1 (.I(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09800__A2 (.I(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09803__S (.I(_03970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09801__S (.I(_03970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12892__A1 (.I(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12788__A1 (.I(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10241__I (.I(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09807__I (.I(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11398__A2 (.I(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11082__A2 (.I(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10018__A1 (.I(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09808__A2 (.I(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14139__A1 (.I(_03980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13526__A1 (.I(_03980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11144__A2 (.I(_03980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09815__A2 (.I(_03980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09818__S (.I(_03981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09816__S (.I(_03981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11903__I (.I(_03984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11058__I (.I(_03984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09821__I (.I(_03984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12899__A1 (.I(_03985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12801__A1 (.I(_03985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10254__I (.I(_03985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09822__I (.I(_03985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13115__A2 (.I(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11205__A2 (.I(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10029__A1 (.I(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09823__A2 (.I(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09826__S (.I(_03987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09824__S (.I(_03987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10665__A1 (.I(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10468__A1 (.I(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10040__A1 (.I(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09835__A1 (.I(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11840__A1 (.I(_03993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11468__A1 (.I(_03993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10662__A1 (.I(_03993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09832__A2 (.I(_03993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09842__I (.I(_03994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09833__I (.I(_03994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10012__I (.I(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09967__I (.I(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09887__I (.I(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09834__I (.I(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11963__A2 (.I(_03996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09877__A1 (.I(_03996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09849__A2 (.I(_03996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09835__A2 (.I(_03996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09857__I0 (.I(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09852__I0 (.I(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09847__I0 (.I(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09839__I0 (.I(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09869__I0 (.I(_04001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09862__I0 (.I(_04001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09855__I0 (.I(_04001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09845__I0 (.I(_04001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10024__A2 (.I(_04002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09930__I (.I(_04002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09894__I (.I(_04002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09843__I (.I(_04002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10055__A1 (.I(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09986__A1 (.I(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09925__A1 (.I(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09861__A1 (.I(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12347__A1 (.I(_04014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11848__A1 (.I(_04014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11133__A1 (.I(_04014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09861__A2 (.I(_04014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09885__I0 (.I(_04018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09880__I0 (.I(_04018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09871__I0 (.I(_04018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09866__I0 (.I(_04018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09871__S (.I(_04020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09869__S (.I(_04020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09908__I0 (.I(_04023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09896__I0 (.I(_04023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09883__I0 (.I(_04023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09878__I0 (.I(_04023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12607__I (.I(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11107__I (.I(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09875__I (.I(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14217__A1 (.I(_04025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11968__A1 (.I(_04025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10077__I (.I(_04025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09876__I (.I(_04025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12011__A2 (.I(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11992__A2 (.I(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11642__A2 (.I(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09877__A2 (.I(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09880__S (.I(_04027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09878__S (.I(_04027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09885__S (.I(_04030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09883__S (.I(_04030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12474__A2 (.I(_04033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09939__A1 (.I(_04033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09900__A2 (.I(_04033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09888__A2 (.I(_04033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09892__S (.I(_04034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09890__A2 (.I(_04034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09889__A2 (.I(_04034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09910__I0 (.I(_04036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09905__I0 (.I(_04036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09898__I0 (.I(_04036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09892__I0 (.I(_04036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09920__A2 (.I(_04038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09914__A2 (.I(_04038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09907__A2 (.I(_04038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09895__A2 (.I(_04038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10469__I (.I(_04043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10281__I (.I(_04043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10108__I (.I(_04043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09902__I (.I(_04043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10093__A1 (.I(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10041__A1 (.I(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09940__A1 (.I(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09903__A1 (.I(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10011__I (.I(_04050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09980__I (.I(_04050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09945__I (.I(_04050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09913__I (.I(_04050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09932__I0 (.I(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09926__I0 (.I(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09921__I0 (.I(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09915__I0 (.I(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09918__S (.I(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09915__S (.I(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09934__I0 (.I(_04054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09928__I0 (.I(_04054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09923__I0 (.I(_04054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09918__I0 (.I(_04054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09934__S (.I(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09932__S (.I(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13924__A1 (.I(_04067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13047__A1 (.I(_04067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11167__I (.I(_04067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09938__I (.I(_04067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11987__A2 (.I(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10261__A2 (.I(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10147__A1 (.I(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09939__A2 (.I(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09965__I0 (.I(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09960__I0 (.I(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09949__I0 (.I(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09943__I0 (.I(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09969__I0 (.I(_04073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09963__I0 (.I(_04073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09958__I0 (.I(_04073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09947__I0 (.I(_04073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09999__A1 (.I(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09975__A2 (.I(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09952__A2 (.I(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10068__I (.I(_04090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10043__I (.I(_04090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10008__I (.I(_04090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09972__I (.I(_04090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09994__I0 (.I(_04091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09989__I0 (.I(_04091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09984__I0 (.I(_04091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09973__I0 (.I(_04091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09978__S (.I(_04093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09976__S (.I(_04093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10006__I0 (.I(_04096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09992__I0 (.I(_04096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09987__I0 (.I(_04096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09982__I0 (.I(_04096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09989__S (.I(_04100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09987__S (.I(_04100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13105__A1 (.I(_04107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13059__A1 (.I(_04107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11229__I (.I(_04107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09998__I (.I(_04107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11974__A2 (.I(_04108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10888__A2 (.I(_04108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10223__A1 (.I(_04108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09999__A2 (.I(_04108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10003__S (.I(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10001__A2 (.I(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10000__A2 (.I(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10226__I1 (.I(_04111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10171__I1 (.I(_04111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10027__I1 (.I(_04111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10003__I1 (.I(_04111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10049__I0 (.I(_04117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10030__I0 (.I(_04117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10019__I0 (.I(_04117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10014__I0 (.I(_04117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10016__S (.I(_04119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10014__S (.I(_04119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10021__S (.I(_04122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10019__S (.I(_04122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12209__A2 (.I(_04125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11255__I (.I(_04125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10247__I (.I(_04125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10024__A1 (.I(_04125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10027__S (.I(_04126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10025__S (.I(_04126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10032__S (.I(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10030__S (.I(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10662__A2 (.I(_04132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10465__A2 (.I(_04132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10269__A1 (.I(_04132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10037__A2 (.I(_04132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10268__A2 (.I(_04133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10036__I (.I(_04133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10046__I (.I(_04135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10038__I (.I(_04135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10215__I (.I(_04136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10174__I (.I(_04136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10091__I (.I(_04136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10039__I (.I(_04136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12369__A2 (.I(_04137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10255__A2 (.I(_04137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10248__A2 (.I(_04137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10040__A2 (.I(_04137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10063__I0 (.I(_04140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10058__I0 (.I(_04140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10051__I0 (.I(_04140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10044__I0 (.I(_04140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12391__A2 (.I(_04142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10130__I (.I(_04142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10078__I (.I(_04142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10047__I (.I(_04142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10071__A2 (.I(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10065__A2 (.I(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10060__A2 (.I(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10048__A2 (.I(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10072__I0 (.I(_04148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10066__I0 (.I(_04148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10061__I0 (.I(_04148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10056__I0 (.I(_04148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10058__S (.I(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10056__S (.I(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10088__I0 (.I(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10082__I0 (.I(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10074__I0 (.I(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10069__I0 (.I(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10115__I0 (.I(_04162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10102__I0 (.I(_04162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10086__I0 (.I(_04162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10080__I0 (.I(_04162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10899__A1 (.I(_04163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10507__A1 (.I(_04163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10306__A1 (.I(_04163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10079__A1 (.I(_04163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10082__S (.I(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10080__S (.I(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10708__A1 (.I(_04168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10514__A1 (.I(_04168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10312__A1 (.I(_04168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10085__A1 (.I(_04168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10088__S (.I(_04169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10086__S (.I(_04169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10911__A1 (.I(_04172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10713__A1 (.I(_04172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10318__A1 (.I(_04172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10092__A1 (.I(_04172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10098__S (.I(_04174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10094__A2 (.I(_04174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10093__A2 (.I(_04174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10456__I (.I(_04176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10331__I (.I(_04176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10219__I (.I(_04176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10096__I (.I(_04176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10117__I0 (.I(_04178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10111__I0 (.I(_04178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10104__I0 (.I(_04178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10098__I0 (.I(_04178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10718__A1 (.I(_04180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10524__A1 (.I(_04180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10323__A1 (.I(_04180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10101__A1 (.I(_04180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10923__A1 (.I(_04184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10724__A1 (.I(_04184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10529__A1 (.I(_04184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10107__A1 (.I(_04184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10111__S (.I(_04185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10110__A2 (.I(_04185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10109__A2 (.I(_04185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10730__A1 (.I(_04189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10535__A1 (.I(_04189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10337__A1 (.I(_04189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10114__A1 (.I(_04189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10143__I0 (.I(_04193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10137__I0 (.I(_04193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10132__I0 (.I(_04193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10124__I0 (.I(_04193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11268__I (.I(_04194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10121__I (.I(_04194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11398__A1 (.I(_04196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11335__A1 (.I(_04196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10760__A1 (.I(_04196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10123__A1 (.I(_04196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10145__I0 (.I(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10139__I0 (.I(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10134__I0 (.I(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10127__I0 (.I(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10744__A1 (.I(_04201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10547__A1 (.I(_04201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10349__A1 (.I(_04201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10131__A1 (.I(_04201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10155__A2 (.I(_04202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10142__A2 (.I(_04202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10136__A2 (.I(_04202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10131__A2 (.I(_04202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10755__A1 (.I(_04209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10560__A1 (.I(_04209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10362__A1 (.I(_04209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10142__A1 (.I(_04209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10184__I0 (.I(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10178__I0 (.I(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10158__I0 (.I(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10151__I0 (.I(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10188__I0 (.I(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10182__I0 (.I(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10176__I0 (.I(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10156__I0 (.I(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10766__A1 (.I(_04218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10572__A1 (.I(_04218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10374__A1 (.I(_04218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10155__A1 (.I(_04218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13406__A1 (.I(_04223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11839__A2 (.I(_04223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10973__A2 (.I(_04223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10163__A1 (.I(_04223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10774__A2 (.I(_04225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10602__A2 (.I(_04225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10382__A1 (.I(_04225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10166__A1 (.I(_04225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12219__A2 (.I(_04226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11667__A1 (.I(_04226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10165__I (.I(_04226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12234__A2 (.I(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11764__A1 (.I(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10974__A1 (.I(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10166__A2 (.I(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12415__A2 (.I(_04228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10223__A2 (.I(_04228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10167__A2 (.I(_04228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10171__S (.I(_04229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10170__A2 (.I(_04229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10169__A2 (.I(_04229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10397__A1 (.I(_04230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10384__A1 (.I(_04230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10224__A1 (.I(_04230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10169__A1 (.I(_04230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10781__A1 (.I(_04233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10584__A1 (.I(_04233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10389__A1 (.I(_04233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10175__A1 (.I(_04233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10987__A1 (.I(_04238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10786__A1 (.I(_04238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10589__A1 (.I(_04238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10181__A1 (.I(_04238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10184__S (.I(_04239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10182__S (.I(_04239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10791__A1 (.I(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10596__A1 (.I(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10401__A1 (.I(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10187__A1 (.I(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10212__I0 (.I(_04245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10207__I0 (.I(_04245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10201__I0 (.I(_04245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10191__I0 (.I(_04245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10594__I (.I(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10488__I (.I(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10335__I (.I(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10194__I (.I(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10304__I (.I(_04248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10266__I (.I(_04248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10234__I (.I(_04248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10195__I (.I(_04248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10230__I0 (.I(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10217__I0 (.I(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10205__I0 (.I(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10199__I0 (.I(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11014__I (.I(_04250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10577__I (.I(_04250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10260__I (.I(_04250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10197__I (.I(_04250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10519__A1 (.I(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10453__A1 (.I(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10328__A1 (.I(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10198__A1 (.I(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10201__S (.I(_04252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10199__S (.I(_04252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10804__A1 (.I(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10611__A1 (.I(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10413__A1 (.I(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10204__A1 (.I(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10207__S (.I(_04256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10205__S (.I(_04256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10817__A1 (.I(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10625__A1 (.I(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10424__A1 (.I(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10216__A1 (.I(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10242__A2 (.I(_04263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10236__A2 (.I(_04263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10229__A2 (.I(_04263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10216__A2 (.I(_04263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10245__I0 (.I(_04267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10239__I0 (.I(_04267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10232__I0 (.I(_04267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10221__I0 (.I(_04267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10226__S (.I(_04269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10225__A2 (.I(_04269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10224__A2 (.I(_04269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10828__A1 (.I(_04272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10635__A1 (.I(_04272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10437__A1 (.I(_04272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10229__A1 (.I(_04272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11042__A1 (.I(_04277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10834__A1 (.I(_04277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10442__A1 (.I(_04277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10236__A1 (.I(_04277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10239__S (.I(_04278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10237__S (.I(_04278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10840__A1 (.I(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10646__A1 (.I(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10448__A1 (.I(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10242__A1 (.I(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10245__S (.I(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10243__S (.I(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11053__A1 (.I(_04285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10845__A1 (.I(_04285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10652__A1 (.I(_04285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10248__A1 (.I(_04285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10252__S (.I(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10249__S (.I(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10275__I0 (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10264__I0 (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10258__I0 (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10252__I0 (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10852__A1 (.I(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10657__A1 (.I(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10460__A1 (.I(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10255__A1 (.I(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10258__S (.I(_04291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10256__S (.I(_04291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12068__A1 (.I(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12011__A1 (.I(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11826__A1 (.I(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10261__A1 (.I(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10264__S (.I(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10263__A2 (.I(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10262__A2 (.I(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10300__I0 (.I(_04298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10294__I0 (.I(_04298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10289__I0 (.I(_04298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10273__I0 (.I(_04298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10870__A1 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10672__A1 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10476__A1 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10272__A1 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10278__I (.I(_04301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10270__I (.I(_04301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12525__A2 (.I(_04302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10343__I (.I(_04302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10305__I (.I(_04302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10271__I (.I(_04302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10876__A1 (.I(_04307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10679__A1 (.I(_04307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10482__A1 (.I(_04307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10280__A1 (.I(_04307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10423__I (.I(_04308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10373__I (.I(_04308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10317__I (.I(_04308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10279__I (.I(_04308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10285__S (.I(_04310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10283__A2 (.I(_04310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10282__A2 (.I(_04310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10419__A1 (.I(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10369__A1 (.I(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10319__A1 (.I(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10282__A1 (.I(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10302__I0 (.I(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10296__I0 (.I(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10291__I0 (.I(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10285__I0 (.I(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10881__A1 (.I(_04315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10685__A1 (.I(_04315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10490__A1 (.I(_04315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10288__A1 (.I(_04315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10296__S (.I(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10294__S (.I(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10893__A1 (.I(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10695__A1 (.I(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10501__A1 (.I(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10299__A1 (.I(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10302__S (.I(_04323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10300__S (.I(_04323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10329__I0 (.I(_04326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10324__I0 (.I(_04326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10313__I0 (.I(_04326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10307__I0 (.I(_04326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10310__S (.I(_04328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10307__S (.I(_04328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10326__I0 (.I(_04330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10321__I0 (.I(_04330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10315__I0 (.I(_04330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10310__I0 (.I(_04330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10315__S (.I(_04332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10313__S (.I(_04332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12396__A2 (.I(_04335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10418__A2 (.I(_04335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10368__A2 (.I(_04335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10318__A2 (.I(_04335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10321__S (.I(_04336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10320__A2 (.I(_04336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10319__A2 (.I(_04336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10333__S (.I(_04342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10329__S (.I(_04342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10352__I0 (.I(_04345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10347__I0 (.I(_04345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10340__I0 (.I(_04345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10333__I0 (.I(_04345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10447__I (.I(_04347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10412__I (.I(_04347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10361__I (.I(_04347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10336__I (.I(_04347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10356__I0 (.I(_04348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10350__I0 (.I(_04348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10345__I0 (.I(_04348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10338__I0 (.I(_04348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10936__A1 (.I(_04352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10735__A1 (.I(_04352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10542__A1 (.I(_04352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10344__A1 (.I(_04352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11157__A1 (.I(_04360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10750__A1 (.I(_04360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10552__A1 (.I(_04360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10355__A1 (.I(_04360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10359__S (.I(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10356__S (.I(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10377__I0 (.I(_04363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10371__I0 (.I(_04363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10365__I0 (.I(_04363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10359__I0 (.I(_04363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10402__I0 (.I(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10390__I0 (.I(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10375__I0 (.I(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10363__I0 (.I(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11373__A1 (.I(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10960__A1 (.I(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10565__A1 (.I(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10368__A1 (.I(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11765__A1 (.I(_04377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11385__A1 (.I(_04377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10975__A1 (.I(_04377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10383__A1 (.I(_04377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11860__A2 (.I(_04378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10381__I (.I(_04378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12166__A1 (.I(_04379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12159__A2 (.I(_04379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11180__A1 (.I(_04379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10382__A2 (.I(_04379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10431__A2 (.I(_04380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10407__A2 (.I(_04380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10383__A2 (.I(_04380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10387__S (.I(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10385__A2 (.I(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10384__A2 (.I(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10435__I1 (.I(_04383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10410__I1 (.I(_04383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10399__I1 (.I(_04383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10387__I1 (.I(_04383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10421__I0 (.I(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10416__I0 (.I(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10404__I0 (.I(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10393__I0 (.I(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10888__A1 (.I(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10640__A2 (.I(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10396__A1 (.I(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10399__S (.I(_04390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10398__A2 (.I(_04390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10397__A2 (.I(_04390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10776__I1 (.I(_04396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10641__I1 (.I(_04396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10604__I1 (.I(_04396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10408__I1 (.I(_04396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10410__S (.I(_04397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10408__S (.I(_04397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10443__I0 (.I(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10438__I0 (.I(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10425__I0 (.I(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10414__I0 (.I(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10451__I0 (.I(_04410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10445__I0 (.I(_04410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10440__I0 (.I(_04410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10428__I0 (.I(_04410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11431__A1 (.I(_04412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11026__A1 (.I(_04412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10630__A1 (.I(_04412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10431__A1 (.I(_04412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10435__S (.I(_04413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10434__A2 (.I(_04413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10433__A2 (.I(_04413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10976__A1 (.I(_04414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10889__A1 (.I(_04414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10631__A1 (.I(_04414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10433__A1 (.I(_04414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10477__I0 (.I(_04423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10461__I0 (.I(_04423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10454__I0 (.I(_04423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10449__I0 (.I(_04423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10458__S (.I(_04427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10454__S (.I(_04427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10532__I (.I(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10510__I (.I(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10485__I (.I(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10457__I (.I(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10479__I0 (.I(_04430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10472__I0 (.I(_04430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10463__I0 (.I(_04430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10458__I0 (.I(_04430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10474__I (.I(_04435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10466__I (.I(_04435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12467__A2 (.I(_04437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10657__A2 (.I(_04437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10652__A2 (.I(_04437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10468__A2 (.I(_04437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10566__A1 (.I(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10530__A1 (.I(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10483__A1 (.I(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10470__A1 (.I(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12427__A2 (.I(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10541__I (.I(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10506__I (.I(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10475__I (.I(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10618__A2 (.I(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10565__A2 (.I(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10529__A2 (.I(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10482__A2 (.I(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10508__I0 (.I(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10502__I0 (.I(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10497__I0 (.I(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10491__I0 (.I(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11298__A1 (.I(_04457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11095__A1 (.I(_04457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10690__A1 (.I(_04457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10496__A1 (.I(_04457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10527__I0 (.I(_04467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10522__I0 (.I(_04467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10517__I0 (.I(_04467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10511__I0 (.I(_04467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10536__I0 (.I(_04469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10525__I0 (.I(_04469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10520__I0 (.I(_04469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10515__I0 (.I(_04469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10522__S (.I(_04473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10520__S (.I(_04473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10550__I0 (.I(_04481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10545__I0 (.I(_04481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10538__I0 (.I(_04481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10533__I0 (.I(_04481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10884__I (.I(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10769__I (.I(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10675__I (.I(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10556__I (.I(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10575__I0 (.I(_04498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10568__I0 (.I(_04498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10563__I0 (.I(_04498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10558__I0 (.I(_04498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10590__I0 (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10585__I0 (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10579__I0 (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10573__I0 (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10596__A2 (.I(_04507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10589__A2 (.I(_04507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10584__A2 (.I(_04507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10572__A2 (.I(_04507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10582__S (.I(_04512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10579__S (.I(_04512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10599__I0 (.I(_04514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10592__I0 (.I(_04514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10587__I0 (.I(_04514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10582__I0 (.I(_04514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10706__I (.I(_04522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10684__I (.I(_04522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10645__I (.I(_04522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10595__I (.I(_04522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10636__I0 (.I(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10626__I0 (.I(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10612__I0 (.I(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10597__I0 (.I(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11001__A1 (.I(_04527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10797__A1 (.I(_04527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10640__A1 (.I(_04527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10603__A1 (.I(_04527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12531__A2 (.I(_04528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10630__A2 (.I(_04528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10603__A2 (.I(_04528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10608__S (.I(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10604__S (.I(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11388__I (.I(_04531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11030__I (.I(_04531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10800__I (.I(_04531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10607__I (.I(_04531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10778__I1 (.I(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10643__I1 (.I(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10633__I1 (.I(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10608__I1 (.I(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10646__A2 (.I(_04534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10635__A2 (.I(_04534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10625__A2 (.I(_04534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10611__A2 (.I(_04534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10638__I0 (.I(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10628__I0 (.I(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10623__I0 (.I(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10615__I0 (.I(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11803__A1 (.I(_04539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11616__A1 (.I(_04539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11419__A1 (.I(_04539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10618__A1 (.I(_04539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11324__I (.I(_04541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10924__I (.I(_04541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10725__I (.I(_04541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10620__I (.I(_04541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10714__A1 (.I(_04542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10680__A1 (.I(_04542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10666__A1 (.I(_04542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10621__A1 (.I(_04542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10633__S (.I(_04548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10632__A2 (.I(_04548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10631__A2 (.I(_04548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10673__I0 (.I(_04557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10658__I0 (.I(_04557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10653__I0 (.I(_04557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10647__I0 (.I(_04557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10668__I0 (.I(_04560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10660__I0 (.I(_04560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10655__I0 (.I(_04560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10650__I0 (.I(_04560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10670__I (.I(_04568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10663__I (.I(_04568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12910__A2 (.I(_04570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10713__A2 (.I(_04570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10679__A2 (.I(_04570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10665__A2 (.I(_04570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10668__S (.I(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10667__A2 (.I(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10666__A2 (.I(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10743__I (.I(_04574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10724__A2 (.I(_04574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10707__I (.I(_04574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10671__I (.I(_04574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10695__A2 (.I(_04575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10690__A2 (.I(_04575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10685__A2 (.I(_04575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10672__A2 (.I(_04575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10747__I (.I(_04578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10721__I (.I(_04578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10698__I (.I(_04578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10676__I (.I(_04578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10693__I0 (.I(_04579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10688__I0 (.I(_04579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10682__I0 (.I(_04579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10677__I0 (.I(_04579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10702__I0 (.I(_04584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10696__I0 (.I(_04584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10691__I0 (.I(_04584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10686__I0 (.I(_04584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10716__I0 (.I(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10711__I0 (.I(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10704__I0 (.I(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10699__I0 (.I(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10704__S (.I(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10702__S (.I(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10736__I0 (.I(_04598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10731__I0 (.I(_04598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10719__I0 (.I(_04598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10709__I0 (.I(_04598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10735__A2 (.I(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10730__A2 (.I(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10718__A2 (.I(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10708__A2 (.I(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10738__I0 (.I(_04608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10733__I0 (.I(_04608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10728__I0 (.I(_04608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10722__I0 (.I(_04608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10912__A1 (.I(_04611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10877__A1 (.I(_04611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10864__A1 (.I(_04611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10726__A1 (.I(_04611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11120__I (.I(_04620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11006__I (.I(_04620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10850__I (.I(_04620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10741__I (.I(_04620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10827__I (.I(_04621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10803__I (.I(_04621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10765__I (.I(_04621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10742__I (.I(_04621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10761__I0 (.I(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10756__I0 (.I(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10751__I0 (.I(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10745__I0 (.I(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10766__A2 (.I(_04623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10755__A2 (.I(_04623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10750__A2 (.I(_04623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10744__A2 (.I(_04623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10763__I0 (.I(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10758__I0 (.I(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10753__I0 (.I(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10748__I0 (.I(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10792__I0 (.I(_04637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10787__I0 (.I(_04637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10782__I0 (.I(_04637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10767__I0 (.I(_04637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10771__S (.I(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10767__S (.I(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10855__I (.I(_04640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10831__I (.I(_04640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10807__I (.I(_04640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10770__I (.I(_04640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10794__I0 (.I(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10789__I0 (.I(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10784__I0 (.I(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10771__I0 (.I(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12702__A2 (.I(_04643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12692__A1 (.I(_04643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11181__A1 (.I(_04643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10775__A1 (.I(_04643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12915__A2 (.I(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10797__A2 (.I(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10775__A2 (.I(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10778__S (.I(_04645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10776__S (.I(_04645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11182__I1 (.I(_04658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11145__I1 (.I(_04658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11002__I1 (.I(_04658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10798__I1 (.I(_04658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10801__S (.I(_04659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10798__S (.I(_04659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11004__I1 (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10978__I1 (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10891__I1 (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10801__I1 (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10823__I0 (.I(_04663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10818__I0 (.I(_04663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10813__I0 (.I(_04663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10805__I0 (.I(_04663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10825__I0 (.I(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10820__I0 (.I(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10815__I0 (.I(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10808__I0 (.I(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12759__A1 (.I(_04668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12709__A2 (.I(_04668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11216__A1 (.I(_04668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10812__A1 (.I(_04668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10834__A2 (.I(_04669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10828__A2 (.I(_04669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10817__A2 (.I(_04669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10812__A2 (.I(_04669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10848__I0 (.I(_04682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10843__I0 (.I(_04682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10837__I0 (.I(_04682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10832__I0 (.I(_04682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12868__A2 (.I(_04687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10852__A2 (.I(_04687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10845__A2 (.I(_04687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10840__A2 (.I(_04687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10843__S (.I(_04688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10841__S (.I(_04688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10894__I0 (.I(_04695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10882__I0 (.I(_04695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10871__I0 (.I(_04695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10853__I0 (.I(_04695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10879__I0 (.I(_04698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10873__I0 (.I(_04698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10866__I0 (.I(_04698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10856__I0 (.I(_04698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12396__A1 (.I(_04700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11682__A1 (.I(_04700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11471__A1 (.I(_04700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10863__A1 (.I(_04700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12928__A2 (.I(_04704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12920__A2 (.I(_04704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11059__A2 (.I(_04704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10863__A2 (.I(_04704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13120__A2 (.I(_04708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10943__I (.I(_04708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10905__I (.I(_04708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10869__I (.I(_04708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10899__A2 (.I(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10893__A2 (.I(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10881__A2 (.I(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10870__A2 (.I(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10960__A2 (.I(_04713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10923__A2 (.I(_04713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10911__A2 (.I(_04713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10876__A2 (.I(_04713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10963__I (.I(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10939__I (.I(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10914__I (.I(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10885__I (.I(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10891__S (.I(_04722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10890__A2 (.I(_04722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10889__A2 (.I(_04722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10931__I0 (.I(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10919__I0 (.I(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10907__I0 (.I(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10900__I0 (.I(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11517__A1 (.I(_04732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11316__A1 (.I(_04732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11113__A1 (.I(_04732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10906__A1 (.I(_04732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11528__A1 (.I(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11329__A1 (.I(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11128__A1 (.I(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10918__A1 (.I(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11288__A1 (.I(_04746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11272__A1 (.I(_04746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10961__A1 (.I(_04746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10925__A1 (.I(_04746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11540__A1 (.I(_04749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11342__A1 (.I(_04749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11138__A1 (.I(_04749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10930__A1 (.I(_04749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10956__I0 (.I(_04753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10950__I0 (.I(_04753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10945__I0 (.I(_04753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10937__I0 (.I(_04753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10940__S (.I(_04754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10937__S (.I(_04754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10958__I0 (.I(_04756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10952__I0 (.I(_04756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10947__I0 (.I(_04756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10940__I0 (.I(_04756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11551__A1 (.I(_04758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11354__A1 (.I(_04758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11150__A1 (.I(_04758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10944__A1 (.I(_04758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10981__A2 (.I(_04759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10968__A2 (.I(_04759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10955__A2 (.I(_04759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10944__A2 (.I(_04759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10947__S (.I(_04760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10945__S (.I(_04760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11564__A1 (.I(_04766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11368__A1 (.I(_04766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11162__A1 (.I(_04766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10955__A1 (.I(_04766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10958__S (.I(_04767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10956__S (.I(_04767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10990__I0 (.I(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10984__I0 (.I(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10971__I0 (.I(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10964__I0 (.I(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10994__I0 (.I(_04774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10988__I0 (.I(_04774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10982__I0 (.I(_04774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10969__I0 (.I(_04774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11576__A1 (.I(_04775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11379__A1 (.I(_04775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11175__A1 (.I(_04775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10968__A1 (.I(_04775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11604__A2 (.I(_04779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11384__A2 (.I(_04779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11180__A2 (.I(_04779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10974__A2 (.I(_04779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11026__A2 (.I(_04780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11001__A2 (.I(_04780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10975__A2 (.I(_04780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11588__A1 (.I(_04784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11391__A1 (.I(_04784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11187__A1 (.I(_04784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10981__A1 (.I(_04784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11598__A1 (.I(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11403__A1 (.I(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11198__A1 (.I(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10993__A1 (.I(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11338__I (.I(_04795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11224__I (.I(_04795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11116__I (.I(_04795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10997__I (.I(_04795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11024__I0 (.I(_04797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11018__I0 (.I(_04797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11012__I0 (.I(_04797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10999__I0 (.I(_04797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11004__S (.I(_04799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11002__S (.I(_04799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11094__I (.I(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11065__I (.I(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11041__I (.I(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11007__I (.I(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11036__I0 (.I(_04803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11022__I0 (.I(_04803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11016__I0 (.I(_04803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11010__I0 (.I(_04803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11611__A1 (.I(_04804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11414__A1 (.I(_04804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11210__A1 (.I(_04804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11009__A1 (.I(_04804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11810__A1 (.I(_04808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11205__A1 (.I(_04808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11082__A1 (.I(_04808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11015__A1 (.I(_04808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11018__S (.I(_04809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11016__S (.I(_04809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11623__A1 (.I(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11426__A1 (.I(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11221__A1 (.I(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11021__A1 (.I(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11630__A1 (.I(_04817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11432__A1 (.I(_04817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11386__A1 (.I(_04817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11028__A1 (.I(_04817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11233__I1 (.I(_04819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11184__I1 (.I(_04819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11147__I1 (.I(_04819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11031__I1 (.I(_04819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11636__A1 (.I(_04821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11437__A1 (.I(_04821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11238__A1 (.I(_04821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11035__A1 (.I(_04821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11053__A2 (.I(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11048__A2 (.I(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11042__A2 (.I(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11035__A2 (.I(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11056__I0 (.I(_04825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11051__I0 (.I(_04825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11045__I0 (.I(_04825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11039__I0 (.I(_04825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11045__S (.I(_04828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11043__S (.I(_04828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11654__A1 (.I(_04831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11447__A1 (.I(_04831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11250__A1 (.I(_04831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11048__A1 (.I(_04831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11675__A1 (.I(_04838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11463__A1 (.I(_04838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11263__A1 (.I(_04838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11059__A1 (.I(_04838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11063__S (.I(_04839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11060__S (.I(_04839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11085__I0 (.I(_04841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11080__I0 (.I(_04841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11074__I0 (.I(_04841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11063__I0 (.I(_04841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11089__I0 (.I(_04843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11083__I0 (.I(_04843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11078__I0 (.I(_04843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11072__I0 (.I(_04843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13615__A1 (.I(_04844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12812__A1 (.I(_04844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11270__I (.I(_04844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11067__I (.I(_04844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12068__A2 (.I(_04845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11912__A1 (.I(_04845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11843__A1 (.I(_04845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11071__A1 (.I(_04845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13417__A2 (.I(_04847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11127__I (.I(_04847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11101__I (.I(_04847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11070__I (.I(_04847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11695__A1 (.I(_04852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11478__A1 (.I(_04852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11279__A1 (.I(_04852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11077__A1 (.I(_04852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11085__S (.I(_04856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11083__S (.I(_04856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11700__A1 (.I(_04859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11492__A1 (.I(_04859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11293__A1 (.I(_04859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11088__A1 (.I(_04859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11092__S (.I(_04860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11089__S (.I(_04860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11111__I0 (.I(_04862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11105__I0 (.I(_04862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11098__I0 (.I(_04862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11092__I0 (.I(_04862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11098__S (.I(_04865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11096__S (.I(_04865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11670__A1 (.I(_04868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11505__A1 (.I(_04868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11304__A1 (.I(_04868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11102__A1 (.I(_04868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11105__S (.I(_04870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11103__S (.I(_04870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12308__A1 (.I(_04873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11512__A1 (.I(_04873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11310__A1 (.I(_04873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11108__A1 (.I(_04873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11111__S (.I(_04874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11109__S (.I(_04874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11118__S (.I(_04877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11114__S (.I(_04877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11201__I (.I(_04879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11171__I (.I(_04879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11141__I (.I(_04879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11117__I (.I(_04879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11136__I0 (.I(_04880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11131__I0 (.I(_04880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11125__I0 (.I(_04880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11118__I0 (.I(_04880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11204__I (.I(_04882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11174__I (.I(_04882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11149__I (.I(_04882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11121__I (.I(_04882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11125__S (.I(_04884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11123__S (.I(_04884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11131__S (.I(_04888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11129__S (.I(_04888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11136__S (.I(_04891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11134__S (.I(_04891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11165__I0 (.I(_04896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11160__I0 (.I(_04896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11153__I0 (.I(_04896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11142__I0 (.I(_04896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11147__S (.I(_04898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11145__S (.I(_04898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11169__I0 (.I(_04901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11163__I0 (.I(_04901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11158__I0 (.I(_04901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11151__I0 (.I(_04901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11153__S (.I(_04902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11151__S (.I(_04902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11249__I (.I(_04905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11215__I (.I(_04905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11186__I (.I(_04905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11156__I (.I(_04905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11175__A2 (.I(_04906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11168__A2 (.I(_04906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11162__A2 (.I(_04906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11157__A2 (.I(_04906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12910__A1 (.I(_04913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12674__A1 (.I(_04913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12570__A2 (.I(_04913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11168__A1 (.I(_04913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11196__I0 (.I(_04916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11190__I0 (.I(_04916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11178__I0 (.I(_04916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11172__I0 (.I(_04916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11199__I0 (.I(_04918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11194__I0 (.I(_04918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11188__I0 (.I(_04918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11176__I0 (.I(_04918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11178__S (.I(_04919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11176__S (.I(_04919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11184__S (.I(_04923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11182__S (.I(_04923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12141__A1 (.I(_04930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11779__A1 (.I(_04930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11593__A1 (.I(_04930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11193__A1 (.I(_04930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11219__I0 (.I(_04936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11213__I0 (.I(_04936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11208__I0 (.I(_04936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11202__I0 (.I(_04936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11222__I0 (.I(_04938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11217__I0 (.I(_04938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11211__I0 (.I(_04938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11206__I0 (.I(_04938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11208__S (.I(_04939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11206__S (.I(_04939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11313__I (.I(_04951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11290__I (.I(_04951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11259__I (.I(_04951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11225__I (.I(_04951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11253__I0 (.I(_04952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11247__I0 (.I(_04952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11241__I0 (.I(_04952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11226__I0 (.I(_04952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11792__I1 (.I(_04954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11606__I1 (.I(_04954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11410__I1 (.I(_04954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11231__I1 (.I(_04954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12915__A1 (.I(_04955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12770__A1 (.I(_04955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12034__A2 (.I(_04955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11230__A1 (.I(_04955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11233__S (.I(_04956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11231__S (.I(_04956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11621__I (.I(_04959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11503__I (.I(_04959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11359__I (.I(_04959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11236__I (.I(_04959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11257__I0 (.I(_04961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11251__I0 (.I(_04961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11245__I0 (.I(_04961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11239__I0 (.I(_04961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12097__A1 (.I(_04965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11882__A1 (.I(_04965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11442__A1 (.I(_04965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11244__A1 (.I(_04965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11247__S (.I(_04966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11245__S (.I(_04966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13164__A2 (.I(_04969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11263__A2 (.I(_04969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11256__A2 (.I(_04969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11250__A2 (.I(_04969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12086__A1 (.I(_04973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11898__A1 (.I(_04973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11659__A1 (.I(_04973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11256__A1 (.I(_04973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11282__I0 (.I(_04976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11274__I0 (.I(_04976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11266__I0 (.I(_04976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11260__I0 (.I(_04976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11299__I0 (.I(_04978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11294__I0 (.I(_04978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11280__I0 (.I(_04978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11264__I0 (.I(_04978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12063__A1 (.I(_04983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11945__A1 (.I(_04983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11744__A1 (.I(_04983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11271__A1 (.I(_04983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13252__A1 (.I(_04984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12275__A1 (.I(_04984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12004__A2 (.I(_04984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11271__A2 (.I(_04984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11285__I (.I(_04988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11277__I (.I(_04988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13620__A2 (.I(_04989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11348__I (.I(_04989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11309__I (.I(_04989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11278__I (.I(_04989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11926__A1 (.I(_04994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11706__A1 (.I(_04994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11485__A1 (.I(_04994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11287__A1 (.I(_04994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11425__I (.I(_04995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11378__I (.I(_04995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11322__I (.I(_04995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11286__I (.I(_04995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14139__A2 (.I(_04996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14077__A2 (.I(_04996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11463__A2 (.I(_04996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11287__A2 (.I(_04996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11291__S (.I(_04997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11289__A2 (.I(_04997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11288__A2 (.I(_04997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11307__I0 (.I(_04999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11301__I0 (.I(_04999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11296__I0 (.I(_04999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11291__I0 (.I(_04999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11330__I0 (.I(_05007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11317__I0 (.I(_05007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11311__I0 (.I(_05007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11305__I0 (.I(_05007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11332__I0 (.I(_05014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11327__I0 (.I(_05014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11319__I0 (.I(_05014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11314__I0 (.I(_05014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12427__A1 (.I(_05019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12222__A1 (.I(_05019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11997__A1 (.I(_05019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11323__A1 (.I(_05019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11327__S (.I(_05021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11326__A2 (.I(_05021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11325__A2 (.I(_05021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11472__A1 (.I(_05022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11420__A1 (.I(_05022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11374__A1 (.I(_05022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11325__A1 (.I(_05022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11355__I0 (.I(_05028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11350__I0 (.I(_05028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11343__I0 (.I(_05028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11336__I0 (.I(_05028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11422__I (.I(_05031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11394__I (.I(_05031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11365__I (.I(_05031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11339__I (.I(_05031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11357__I0 (.I(_05032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11352__I0 (.I(_05032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11345__I0 (.I(_05032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11340__I0 (.I(_05032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12322__A1 (.I(_05037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11720__A1 (.I(_05037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11546__A1 (.I(_05037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11349__A1 (.I(_05037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11462__I (.I(_05045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11436__I (.I(_05045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11397__I (.I(_05045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11360__I (.I(_05045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11392__I0 (.I(_05046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11380__I0 (.I(_05046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11369__I0 (.I(_05046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11363__I0 (.I(_05046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11958__A1 (.I(_05047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11731__A1 (.I(_05047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11559__A1 (.I(_05047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11362__A1 (.I(_05047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11366__S (.I(_05048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11363__S (.I(_05048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11382__I0 (.I(_05050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11376__I0 (.I(_05050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11371__I0 (.I(_05050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11366__I0 (.I(_05050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11376__S (.I(_05055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11375__A2 (.I(_05055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11374__A2 (.I(_05055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11414__A2 (.I(_05058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11403__A2 (.I(_05058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11391__A2 (.I(_05058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11379__A2 (.I(_05058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11431__A2 (.I(_05062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11409__A2 (.I(_05062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11385__A2 (.I(_05062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11608__I1 (.I(_05065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11434__I1 (.I(_05065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11412__I1 (.I(_05065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11389__I1 (.I(_05065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11417__I0 (.I(_05069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11406__I0 (.I(_05069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11401__I0 (.I(_05069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11395__I0 (.I(_05069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11427__I0 (.I(_05071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11415__I0 (.I(_05071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11404__I0 (.I(_05071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11399__I0 (.I(_05071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11933__A1 (.I(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11791__A1 (.I(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11605__A1 (.I(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11409__A1 (.I(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11423__S (.I(_05085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11421__A2 (.I(_05085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11420__A2 (.I(_05085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11445__I0 (.I(_05087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11440__I0 (.I(_05087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11429__I0 (.I(_05087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11423__I0 (.I(_05087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11458__I0 (.I(_05096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11448__I0 (.I(_05096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11443__I0 (.I(_05096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11438__I0 (.I(_05096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12791__I (.I(_05105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12336__I (.I(_05105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11885__I (.I(_05105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11451__I (.I(_05105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11775__I (.I(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11662__I (.I(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11554__I (.I(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11452__I (.I(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11531__I (.I(_05107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11508__I (.I(_05107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11481__I (.I(_05107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11453__I (.I(_05107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11474__I0 (.I(_05108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11466__I0 (.I(_05108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11460__I0 (.I(_05108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11454__I0 (.I(_05108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11642__A1 (.I(_05110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11582__A1 (.I(_05110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11522__A1 (.I(_05110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11457__A1 (.I(_05110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11460__S (.I(_05111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11458__S (.I(_05111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11499__I0 (.I(_05114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11493__I0 (.I(_05114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11479__I0 (.I(_05114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11464__I0 (.I(_05114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11476__I (.I(_05118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11469__I (.I(_05118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11610__I (.I(_05119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11575__I (.I(_05119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11484__I (.I(_05119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11470__I (.I(_05119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14212__A2 (.I(_05120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11675__A2 (.I(_05120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11659__A2 (.I(_05120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11471__A2 (.I(_05120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14182__A2 (.I(_05124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11545__I (.I(_05124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11511__I (.I(_05124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11477__I (.I(_05124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11501__I0 (.I(_05128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11495__I0 (.I(_05128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11490__I0 (.I(_05128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11482__I0 (.I(_05128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11616__A2 (.I(_05130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11570__A2 (.I(_05130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11535__A2 (.I(_05130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11485__A2 (.I(_05130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11946__I (.I(_05132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11804__I (.I(_05132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11683__I (.I(_05132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11487__I (.I(_05132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11617__A1 (.I(_05133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11571__A1 (.I(_05133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11536__A1 (.I(_05133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11488__A1 (.I(_05133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12297__A1 (.I(_05139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11963__A1 (.I(_05139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11689__A1 (.I(_05139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11498__A1 (.I(_05139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11501__S (.I(_05140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11499__S (.I(_05140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11523__I0 (.I(_05144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11518__I0 (.I(_05144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11513__I0 (.I(_05144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11506__I0 (.I(_05144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11509__S (.I(_05145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11506__S (.I(_05145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11525__I0 (.I(_05147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11520__I0 (.I(_05147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11515__I0 (.I(_05147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11509__I0 (.I(_05147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11515__S (.I(_05150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11513__S (.I(_05150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11520__S (.I(_05153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11518__S (.I(_05153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11525__S (.I(_05156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11523__S (.I(_05156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11552__I0 (.I(_05159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11547__I0 (.I(_05159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11541__I0 (.I(_05159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11529__I0 (.I(_05159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11549__I0 (.I(_05162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11543__I0 (.I(_05162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11538__I0 (.I(_05162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11532__I0 (.I(_05162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13620__A1 (.I(_05164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12525__A1 (.I(_05164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12044__A1 (.I(_05164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11535__A1 (.I(_05164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11573__I0 (.I(_05178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11567__I0 (.I(_05178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11562__I0 (.I(_05178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11556__I0 (.I(_05178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11583__I0 (.I(_05180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11577__I0 (.I(_05180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11565__I0 (.I(_05180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11560__I0 (.I(_05180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11562__S (.I(_05181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11560__S (.I(_05181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11567__S (.I(_05184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11565__S (.I(_05184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12408__A1 (.I(_05187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12146__A1 (.I(_05187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11758__A1 (.I(_05187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11570__A1 (.I(_05187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11573__S (.I(_05188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11572__A2 (.I(_05188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11571__A2 (.I(_05188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11598__A2 (.I(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11593__A2 (.I(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11588__A2 (.I(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11576__A2 (.I(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11580__S (.I(_05192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11577__S (.I(_05192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11596__I0 (.I(_05194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11591__I0 (.I(_05194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11585__I0 (.I(_05194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11580__I0 (.I(_05194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11585__S (.I(_05196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11583__S (.I(_05196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11612__I0 (.I(_05199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11599__I0 (.I(_05199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11594__I0 (.I(_05199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11589__I0 (.I(_05199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11602__S (.I(_05206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11599__S (.I(_05206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11626__I0 (.I(_05208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11619__I0 (.I(_05208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11614__I0 (.I(_05208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11602__I0 (.I(_05208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14207__A2 (.I(_05210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11629__A2 (.I(_05210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11605__A2 (.I(_05210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11608__S (.I(_05211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11606__S (.I(_05211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11614__S (.I(_05215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11612__S (.I(_05215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11719__I (.I(_05221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11688__I (.I(_05221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11653__I (.I(_05221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11622__I (.I(_05221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11649__I0 (.I(_05222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11643__I0 (.I(_05222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11637__I0 (.I(_05222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11624__I0 (.I(_05222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12806__A1 (.I(_05226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12536__A1 (.I(_05226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12229__A1 (.I(_05226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11629__A1 (.I(_05226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12418__I (.I(_05229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12200__I (.I(_05229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11977__I (.I(_05229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11633__I (.I(_05229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11936__I1 (.I(_05230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11794__I1 (.I(_05230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11769__I1 (.I(_05230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11634__I1 (.I(_05230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11657__I0 (.I(_05234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11651__I0 (.I(_05234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11645__I0 (.I(_05234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11640__I0 (.I(_05234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11645__S (.I(_05236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11643__S (.I(_05236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12029__A1 (.I(_05239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11853__A1 (.I(_05239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11821__A1 (.I(_05239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11648__A1 (.I(_05239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11651__S (.I(_05240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11649__S (.I(_05240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11676__I0 (.I(_05243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11671__I0 (.I(_05243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11660__I0 (.I(_05243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11655__I0 (.I(_05243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11741__I (.I(_05249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11716__I (.I(_05249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11692__I (.I(_05249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11663__I (.I(_05249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11686__I0 (.I(_05250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11678__I0 (.I(_05250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11673__I0 (.I(_05250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11664__I0 (.I(_05250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11763__I (.I(_05252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11667__A2 (.I(_05252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11680__I (.I(_05253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11668__I (.I(_05253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14149__A2 (.I(_05254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11737__I (.I(_05254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11712__I (.I(_05254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11669__I (.I(_05254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11678__S (.I(_05259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11676__S (.I(_05259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11881__I (.I(_05262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11785__I (.I(_05262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11705__I (.I(_05262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11681__I (.I(_05262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14217__A2 (.I(_05263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14187__A2 (.I(_05263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12876__A2 (.I(_05263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11682__A2 (.I(_05263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11714__I0 (.I(_05268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11701__I0 (.I(_05268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11696__I0 (.I(_05268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11690__I0 (.I(_05268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11709__I0 (.I(_05271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11703__I0 (.I(_05271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11698__I0 (.I(_05271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11693__I0 (.I(_05271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14088__A2 (.I(_05279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11803__A2 (.I(_05279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11758__A2 (.I(_05279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11706__A2 (.I(_05279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12614__A1 (.I(_05283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12328__A1 (.I(_05283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11982__A1 (.I(_05283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11713__A1 (.I(_05283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11723__S (.I(_05290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11721__S (.I(_05290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12650__A1 (.I(_05293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12379__A1 (.I(_05293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12116__A1 (.I(_05293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11726__A1 (.I(_05293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11729__S (.I(_05294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11727__S (.I(_05294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11734__S (.I(_05297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11732__S (.I(_05297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12660__A1 (.I(_05300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12402__A1 (.I(_05300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12129__A1 (.I(_05300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11738__A1 (.I(_05300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11742__S (.I(_05302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11739__S (.I(_05302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11761__I0 (.I(_05304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11756__I0 (.I(_05304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11747__I0 (.I(_05304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11742__I0 (.I(_05304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11747__S (.I(_05306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11746__A2 (.I(_05306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11745__A2 (.I(_05306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12182__I (.I(_05309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12056__I (.I(_05309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11896__I (.I(_05309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11750__I (.I(_05309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11787__I0 (.I(_05311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11780__I0 (.I(_05311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11773__I0 (.I(_05311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11754__I0 (.I(_05311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12679__A1 (.I(_05312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12422__A1 (.I(_05312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12153__A1 (.I(_05312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11753__A1 (.I(_05312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12691__A2 (.I(_05319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12166__A2 (.I(_05319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11932__A2 (.I(_05319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11764__A2 (.I(_05319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12806__A2 (.I(_05320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11791__A2 (.I(_05320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11765__A2 (.I(_05320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11769__S (.I(_05321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11768__A2 (.I(_05321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11767__A2 (.I(_05321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12230__A1 (.I(_05322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12168__A1 (.I(_05322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11975__A1 (.I(_05322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11767__A1 (.I(_05322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12437__A1 (.I(_05325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12177__A1 (.I(_05325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12172__A1 (.I(_05325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11772__A1 (.I(_05325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11856__I (.I(_05328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11829__I (.I(_05328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11807__I (.I(_05328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11776__I (.I(_05328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11801__I0 (.I(_05329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11789__I0 (.I(_05329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11782__I0 (.I(_05329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11777__I0 (.I(_05329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11782__S (.I(_05331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11780__S (.I(_05331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12491__A1 (.I(_05334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12192__A1 (.I(_05334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12134__A1 (.I(_05334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11786__A1 (.I(_05334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11834__A2 (.I(_05335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11816__A2 (.I(_05335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11798__A2 (.I(_05335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11786__A2 (.I(_05335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11789__S (.I(_05336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11787__S (.I(_05336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11794__S (.I(_05339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11792__S (.I(_05339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11822__I0 (.I(_05342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11817__I0 (.I(_05342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11811__I0 (.I(_05342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11799__I0 (.I(_05342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12509__A1 (.I(_05343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12203__A1 (.I(_05343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11868__A1 (.I(_05343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11798__A1 (.I(_05343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11801__S (.I(_05344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11799__S (.I(_05344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11927__A1 (.I(_05348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11877__A1 (.I(_05348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11827__A1 (.I(_05348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11805__A1 (.I(_05348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11824__I0 (.I(_05350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11819__I0 (.I(_05350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11813__I0 (.I(_05350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11808__I0 (.I(_05350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11813__S (.I(_05352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11811__S (.I(_05352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12520__A1 (.I(_05355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12214__A1 (.I(_05355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11863__A1 (.I(_05355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11816__A1 (.I(_05355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11824__S (.I(_05359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11822__S (.I(_05359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11830__S (.I(_05362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11828__A2 (.I(_05362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11827__A2 (.I(_05362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11851__I0 (.I(_05364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11846__I0 (.I(_05364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11837__I0 (.I(_05364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11830__I0 (.I(_05364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11854__I0 (.I(_05366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11849__I0 (.I(_05366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11844__I0 (.I(_05366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11835__I0 (.I(_05366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12541__A1 (.I(_05367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12242__A1 (.I(_05367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12110__A1 (.I(_05367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11834__A1 (.I(_05367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12272__A2 (.I(_05371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11909__A2 (.I(_05371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11840__A2 (.I(_05371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12642__I (.I(_05372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11841__I (.I(_05372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13526__A2 (.I(_05373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12613__I (.I(_05373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12587__I (.I(_05373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11842__I (.I(_05373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12582__A2 (.I(_05374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12577__A2 (.I(_05374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11848__A2 (.I(_05374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11843__A2 (.I(_05374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11879__I0 (.I(_05383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11871__I0 (.I(_05383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11866__I0 (.I(_05383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11857__I0 (.I(_05383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11892__I0 (.I(_05385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11883__I0 (.I(_05385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11869__I0 (.I(_05385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11864__I0 (.I(_05385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11874__I (.I(_05386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11861__I (.I(_05386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13047__A2 (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12140__I (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12091__I (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11862__I (.I(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12086__A2 (.I(_05388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12073__A2 (.I(_05388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11868__A2 (.I(_05388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11863__A2 (.I(_05388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12748__A1 (.I(_05395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12514__A1 (.I(_05395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12474__A1 (.I(_05395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11876__A1 (.I(_05395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13240__I (.I(_05396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13035__I (.I(_05396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12886__I (.I(_05396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11875__I (.I(_05396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14171__A2 (.I(_05397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14144__A2 (.I(_05397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14110__A2 (.I(_05397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11876__A2 (.I(_05397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11879__S (.I(_05398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11878__A2 (.I(_05398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11877__A2 (.I(_05398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11888__S (.I(_05402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11883__S (.I(_05402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11971__I (.I(_05405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11949__I (.I(_05405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11915__I (.I(_05405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11887__I (.I(_05405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11907__I0 (.I(_05406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11901__I0 (.I(_05406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11894__I0 (.I(_05406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11888__I0 (.I(_05406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12553__A1 (.I(_05408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12254__A1 (.I(_05408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12092__A1 (.I(_05408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11891__A1 (.I(_05408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11894__S (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11892__S (.I(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11920__I0 (.I(_05413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11913__I0 (.I(_05413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11905__I0 (.I(_05413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11899__I0 (.I(_05413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11901__S (.I(_05414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11899__S (.I(_05414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12563__A1 (.I(_05417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12267__A1 (.I(_05417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12073__A1 (.I(_05417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11904__A1 (.I(_05417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11907__S (.I(_05418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11905__S (.I(_05418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11924__I (.I(_05421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11910__I (.I(_05421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12748__A2 (.I(_05422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12128__I (.I(_05422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11981__I (.I(_05422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11911__I (.I(_05422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11953__A2 (.I(_05423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11940__A2 (.I(_05423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11919__A2 (.I(_05423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11912__A2 (.I(_05423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11943__I0 (.I(_05426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11929__I0 (.I(_05426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11922__I0 (.I(_05426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11916__I0 (.I(_05426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12577__A1 (.I(_05428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12280__A1 (.I(_05428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12058__A1 (.I(_05428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11919__A1 (.I(_05428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12248__I (.I(_05432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12191__I (.I(_05432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12104__I (.I(_05432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11925__I (.I(_05432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11929__S (.I(_05434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11928__A2 (.I(_05434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11927__A2 (.I(_05434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12198__I1 (.I(_05437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12161__I1 (.I(_05437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12035__I1 (.I(_05437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11934__I1 (.I(_05437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12536__A2 (.I(_05438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12432__A2 (.I(_05438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11933__A2 (.I(_05438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11936__S (.I(_05439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11934__S (.I(_05439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11964__I0 (.I(_05442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11959__I0 (.I(_05442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11954__I0 (.I(_05442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11941__I0 (.I(_05442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12588__A1 (.I(_05443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12292__A1 (.I(_05443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12039__A1 (.I(_05443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11940__A1 (.I(_05443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11998__A1 (.I(_05448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11988__A1 (.I(_05448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11969__A1 (.I(_05448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11947__A1 (.I(_05448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11966__I0 (.I(_05450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11961__I0 (.I(_05450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11956__I0 (.I(_05450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11950__I0 (.I(_05450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12354__A1 (.I(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12303__A1 (.I(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12023__A1 (.I(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11953__A1 (.I(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11961__S (.I(_05456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11959__S (.I(_05456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11966__S (.I(_05459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11964__S (.I(_05459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11995__I0 (.I(_05464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11990__I0 (.I(_05464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11985__I0 (.I(_05464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11972__I0 (.I(_05464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12170__I1 (.I(_05468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12163__I1 (.I(_05468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12037__I1 (.I(_05468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11978__I1 (.I(_05468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12018__I0 (.I(_05470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12012__I0 (.I(_05470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11993__I0 (.I(_05470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11983__I0 (.I(_05470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12116__A2 (.I(_05471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12080__A2 (.I(_05471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12017__A2 (.I(_05471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11982__A2 (.I(_05471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11990__S (.I(_05475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11989__A2 (.I(_05475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11988__A2 (.I(_05475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12002__S (.I(_05481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11999__A2 (.I(_05481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11998__A2 (.I(_05481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12020__I0 (.I(_05484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12014__I0 (.I(_05484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12009__I0 (.I(_05484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12002__I0 (.I(_05484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12106__A1 (.I(_05488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12064__A1 (.I(_05488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12045__A1 (.I(_05488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12007__A1 (.I(_05488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12876__A1 (.I(_05494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12626__A1 (.I(_05494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12342__A1 (.I(_05494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12017__A1 (.I(_05494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12051__I0 (.I(_05498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12040__I0 (.I(_05498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12030__I0 (.I(_05498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12024__I0 (.I(_05498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12047__I0 (.I(_05501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12042__I0 (.I(_05501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12032__I0 (.I(_05501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12027__I0 (.I(_05501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12037__S (.I(_05506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12035__S (.I(_05506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12042__S (.I(_05509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12040__S (.I(_05509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12047__S (.I(_05512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12046__A2 (.I(_05512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12045__A2 (.I(_05512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13164__A1 (.I(_05515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12582__A1 (.I(_05515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12317__A1 (.I(_05515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12050__A1 (.I(_05515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12054__S (.I(_05516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12051__S (.I(_05516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12071__I0 (.I(_05518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12066__I0 (.I(_05518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12061__I0 (.I(_05518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12054__I0 (.I(_05518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12081__I0 (.I(_05521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12074__I0 (.I(_05521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12069__I0 (.I(_05521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12059__I0 (.I(_05521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12061__S (.I(_05522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12059__S (.I(_05522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12066__S (.I(_05525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12065__A2 (.I(_05525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12064__A2 (.I(_05525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12071__S (.I(_05528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12069__S (.I(_05528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12095__I0 (.I(_05533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12089__I0 (.I(_05533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12083__I0 (.I(_05533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12077__I0 (.I(_05533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13025__A1 (.I(_05535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12636__A1 (.I(_05535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12361__A1 (.I(_05535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12080__A1 (.I(_05535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12111__I0 (.I(_05539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12098__I0 (.I(_05539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12093__I0 (.I(_05539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12087__I0 (.I(_05539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12134__A2 (.I(_05543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12110__A2 (.I(_05543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12097__A2 (.I(_05543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12092__A2 (.I(_05543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12102__S (.I(_05547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12098__S (.I(_05547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12188__I (.I(_05549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12150__I (.I(_05549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12125__I (.I(_05549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12101__I (.I(_05549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12119__I0 (.I(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12113__I0 (.I(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12108__I0 (.I(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12102__I0 (.I(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12743__A2 (.I(_05552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12737__A2 (.I(_05552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12146__A2 (.I(_05552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12105__A2 (.I(_05552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12108__S (.I(_05553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12107__A2 (.I(_05553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12106__A2 (.I(_05553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12135__I0 (.I(_05559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12130__I0 (.I(_05559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12123__I0 (.I(_05559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12117__I0 (.I(_05559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12503__A1 (.I(_05563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12374__A1 (.I(_05563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12285__A1 (.I(_05563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12122__A1 (.I(_05563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12126__S (.I(_05564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12123__S (.I(_05564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12144__I0 (.I(_05566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12137__I0 (.I(_05566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12132__I0 (.I(_05566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12126__I0 (.I(_05566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12185__A2 (.I(_05568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12177__A2 (.I(_05568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12153__A2 (.I(_05568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12129__A2 (.I(_05568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12178__I0 (.I(_05575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12173__I0 (.I(_05575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12154__I0 (.I(_05575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12142__I0 (.I(_05575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12754__A2 (.I(_05576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12726__A2 (.I(_05576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12172__A2 (.I(_05576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12141__A2 (.I(_05576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12397__A1 (.I(_05581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12392__A1 (.I(_05581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12223__A1 (.I(_05581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12148__A1 (.I(_05581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12180__I0 (.I(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12175__I0 (.I(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12156__I0 (.I(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12151__I0 (.I(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12721__A1 (.I(_05588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12415__A1 (.I(_05588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12197__A1 (.I(_05588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12160__A1 (.I(_05588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13059__A2 (.I(_05589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12684__A2 (.I(_05589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12160__A2 (.I(_05589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12163__S (.I(_05590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12161__S (.I(_05590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12531__A1 (.I(_05593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12432__A1 (.I(_05593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12235__A1 (.I(_05593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12167__A1 (.I(_05593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12229__A2 (.I(_05594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12197__A2 (.I(_05594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12167__A2 (.I(_05594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12170__S (.I(_05595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12169__A2 (.I(_05595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12168__A2 (.I(_05595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12291__I (.I(_05604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12266__I (.I(_05604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12241__I (.I(_05604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12183__I (.I(_05604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12215__I0 (.I(_05605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12204__I0 (.I(_05605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12193__I0 (.I(_05605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12186__I0 (.I(_05605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13041__A1 (.I(_05606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12497__A1 (.I(_05606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12486__A1 (.I(_05606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12185__A1 (.I(_05606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12189__S (.I(_05607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12186__S (.I(_05607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12217__I0 (.I(_05609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12206__I0 (.I(_05609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12195__I0 (.I(_05609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12189__I0 (.I(_05609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12242__A2 (.I(_05611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12214__A2 (.I(_05611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12203__A2 (.I(_05611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12192__A2 (.I(_05611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12201__S (.I(_05615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12198__S (.I(_05615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12239__I1 (.I(_05617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12232__I1 (.I(_05617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12212__I1 (.I(_05617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12201__I1 (.I(_05617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12703__I1 (.I(_05622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12693__I1 (.I(_05622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12416__I1 (.I(_05622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12210__I1 (.I(_05622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12352__I (.I(_05629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12220__I (.I(_05629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14132__A2 (.I(_05631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14127__A2 (.I(_05631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14122__A2 (.I(_05631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12222__A2 (.I(_05631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12227__S (.I(_05632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12224__A2 (.I(_05632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12223__A2 (.I(_05632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12311__I (.I(_05634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12288__I (.I(_05634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12263__I (.I(_05634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12226__I (.I(_05634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12257__I0 (.I(_05635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12252__I0 (.I(_05635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12245__I0 (.I(_05635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12227__I0 (.I(_05635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12232__S (.I(_05637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12231__A2 (.I(_05637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12230__A2 (.I(_05637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13105__A2 (.I(_05640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13075__A2 (.I(_05640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12235__A2 (.I(_05640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12239__S (.I(_05641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12238__A2 (.I(_05641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12237__A2 (.I(_05641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12537__A1 (.I(_05642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12532__A1 (.I(_05642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12433__A1 (.I(_05642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12237__A1 (.I(_05642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12783__A1 (.I(_05649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12547__A1 (.I(_05649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12467__A1 (.I(_05649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12249__A1 (.I(_05649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12905__A1 (.I(_05657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12558__A1 (.I(_05657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12481__A1 (.I(_05657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12260__A1 (.I(_05657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12283__I0 (.I(_05660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12278__I0 (.I(_05660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12270__I0 (.I(_05660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12264__I0 (.I(_05660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12286__I0 (.I(_05662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12281__I0 (.I(_05662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12276__I0 (.I(_05662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12268__I0 (.I(_05662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12359__I (.I(_05666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12273__I (.I(_05666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12514__A2 (.I(_05667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12327__I (.I(_05667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12302__I (.I(_05667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12274__I (.I(_05667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12297__A2 (.I(_05668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12292__A2 (.I(_05668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12280__A2 (.I(_05668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12275__A2 (.I(_05668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12306__I0 (.I(_05677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12300__I0 (.I(_05677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12295__I0 (.I(_05677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12289__I0 (.I(_05677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12309__I0 (.I(_05679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12304__I0 (.I(_05679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12298__I0 (.I(_05679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12293__I0 (.I(_05679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12300__S (.I(_05683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12298__S (.I(_05683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12312__S (.I(_05690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12309__S (.I(_05690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12331__I0 (.I(_05692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12325__I0 (.I(_05692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12320__I0 (.I(_05692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12312__I0 (.I(_05692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12707__I (.I(_05694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12593__I (.I(_05694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12479__I (.I(_05694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12315__I (.I(_05694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12334__I0 (.I(_05696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12329__I0 (.I(_05696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12323__I0 (.I(_05696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12318__I0 (.I(_05696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12320__S (.I(_05697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12318__S (.I(_05697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12325__S (.I(_05700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12323__S (.I(_05700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12347__A2 (.I(_05703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12342__A2 (.I(_05703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12333__A2 (.I(_05703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12328__A2 (.I(_05703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12669__I (.I(_05709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12573__I (.I(_05709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12470__I (.I(_05709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12337__I (.I(_05709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12357__I0 (.I(_05711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12350__I0 (.I(_05711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12345__I0 (.I(_05711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12339__I0 (.I(_05711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12362__I0 (.I(_05713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12355__I0 (.I(_05713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12348__I0 (.I(_05713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12343__I0 (.I(_05713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14105__A2 (.I(_05720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12904__I (.I(_05720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12838__I (.I(_05720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12353__I (.I(_05720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12830__A2 (.I(_05721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12819__A2 (.I(_05721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12666__A2 (.I(_05721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12354__A2 (.I(_05721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12508__I (.I(_05725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12421__I (.I(_05725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12407__I (.I(_05725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12360__I (.I(_05725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12402__A2 (.I(_05726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12385__A2 (.I(_05726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12379__A2 (.I(_05726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12361__A2 (.I(_05726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12365__S (.I(_05727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12362__S (.I(_05727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12382__I0 (.I(_05729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12377__I0 (.I(_05729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12372__I0 (.I(_05729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12365__I0 (.I(_05729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12386__I0 (.I(_05731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12380__I0 (.I(_05731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12375__I0 (.I(_05731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12370__I0 (.I(_05731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13417__A1 (.I(_05732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13036__A1 (.I(_05732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12644__A1 (.I(_05732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12369__A1 (.I(_05732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12372__S (.I(_05733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12370__S (.I(_05733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13069__A1 (.I(_05742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12928__A1 (.I(_05742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12655__A1 (.I(_05742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12385__A1 (.I(_05742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12405__I0 (.I(_05745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12399__I0 (.I(_05745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12394__I0 (.I(_05745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12389__I0 (.I(_05745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12468__I0 (.I(_05753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12438__I0 (.I(_05753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12423__I0 (.I(_05753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12403__I0 (.I(_05753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12563__A2 (.I(_05757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12558__A2 (.I(_05757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12553__A2 (.I(_05757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12408__A2 (.I(_05757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12413__S (.I(_05758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12411__A2 (.I(_05758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12410__A2 (.I(_05758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12515__A1 (.I(_05759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12475__A1 (.I(_05759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12428__A1 (.I(_05759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12410__A1 (.I(_05759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12440__I0 (.I(_05761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12430__I0 (.I(_05761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12425__I0 (.I(_05761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12413__I0 (.I(_05761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12419__S (.I(_05763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12416__S (.I(_05763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12539__I1 (.I(_05765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12534__I1 (.I(_05765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12435__I1 (.I(_05765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12419__I1 (.I(_05765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12491__A2 (.I(_05767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12486__A2 (.I(_05767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12437__A2 (.I(_05767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12422__A2 (.I(_05767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12425__S (.I(_05768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12423__S (.I(_05768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12435__S (.I(_05774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12434__A2 (.I(_05774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12433__A2 (.I(_05774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12440__S (.I(_05777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12438__S (.I(_05777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14169__A1 (.I(_05780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12997__B2 (.I(_05780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12990__A1 (.I(_05780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12450__A1 (.I(_05780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13184__A1 (.I(_05783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13180__A1 (.I(_05783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12959__A2 (.I(_05783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12446__I (.I(_05783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13716__I (.I(_05784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13390__A1 (.I(_05784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12943__A1 (.I(_05784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12448__A2 (.I(_05784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13126__I (.I(_05785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12448__B (.I(_05785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12863__I (.I(_05786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12449__I (.I(_05786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13841__A1 (.I(_05787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13695__I (.I(_05787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13259__A1 (.I(_05787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12450__B (.I(_05787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12844__A1 (.I(_05788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12837__A2 (.I(_05788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12451__A2 (.I(_05788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14168__A1 (.I(_05790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13915__A1 (.I(_05790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13832__A1 (.I(_05790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12464__A1 (.I(_05790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13937__I (.I(_05792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12460__A1 (.I(_05792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12460__B1 (.I(_05797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13972__B2 (.I(_05798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12461__A3 (.I(_05798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13938__A1 (.I(_05800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13934__C (.I(_05800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12463__I (.I(_05800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14001__I (.I(_05801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13966__I (.I(_05801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13931__I (.I(_05801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12464__B (.I(_05801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12465__A4 (.I(_05802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14193__A2 (.I(_05803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12844__A2 (.I(_05803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12466__A2 (.I(_05803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12489__I0 (.I(_05807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12484__I0 (.I(_05807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12477__I0 (.I(_05807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12472__I0 (.I(_05807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12498__I0 (.I(_05813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12492__I0 (.I(_05813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12487__I0 (.I(_05813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12482__I0 (.I(_05813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12512__I0 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12506__I0 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12500__I0 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12495__I0 (.I(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12542__I0 (.I(_05827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12521__I0 (.I(_05827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12510__I0 (.I(_05827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12504__I0 (.I(_05827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12547__A2 (.I(_05831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12541__A2 (.I(_05831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12520__A2 (.I(_05831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12509__A2 (.I(_05831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12518__S (.I(_05835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12516__A2 (.I(_05835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12515__A2 (.I(_05835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12544__I0 (.I(_05837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12529__I0 (.I(_05837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12523__I0 (.I(_05837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12518__I0 (.I(_05837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12749__A1 (.I(_05843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12744__A1 (.I(_05843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12738__A1 (.I(_05843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12527__A1 (.I(_05843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12534__S (.I(_05846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12533__A2 (.I(_05846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12532__A2 (.I(_05846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12539__S (.I(_05849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12538__A2 (.I(_05849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12537__A2 (.I(_05849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12564__I0 (.I(_05855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12559__I0 (.I(_05855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12554__I0 (.I(_05855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12548__I0 (.I(_05855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12551__S (.I(_05856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12548__S (.I(_05856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12566__S (.I(_05866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12564__S (.I(_05866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12589__I0 (.I(_05869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12583__I0 (.I(_05869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12578__I0 (.I(_05869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12571__I0 (.I(_05869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12796__A1 (.I(_05870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12709__A1 (.I(_05870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12631__A1 (.I(_05870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12570__A1 (.I(_05870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12647__I (.I(_05873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12623__I (.I(_05873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12599__I (.I(_05873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12574__I (.I(_05873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12591__I0 (.I(_05874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12585__I0 (.I(_05874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12580__I0 (.I(_05874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12575__I0 (.I(_05874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12608__A2 (.I(_05882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12602__A2 (.I(_05882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12596__A2 (.I(_05882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12588__A2 (.I(_05882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12591__S (.I(_05883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12589__S (.I(_05883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12665__I (.I(_05886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12641__I (.I(_05886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12619__I (.I(_05886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12594__I (.I(_05886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13093__A1 (.I(_05888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12920__A1 (.I(_05888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12839__A1 (.I(_05888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12596__A1 (.I(_05888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12600__S (.I(_05889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12597__S (.I(_05889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12605__S (.I(_05893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12603__S (.I(_05893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12887__A1 (.I(_05896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12868__A1 (.I(_05896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12666__A1 (.I(_05896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12608__A1 (.I(_05896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12611__S (.I(_05897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12609__S (.I(_05897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12617__S (.I(_05901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12615__S (.I(_05901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12637__I0 (.I(_05904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12632__I0 (.I(_05904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12627__I0 (.I(_05904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12621__I0 (.I(_05904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12639__I0 (.I(_05907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12634__I0 (.I(_05907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12629__I0 (.I(_05907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12624__I0 (.I(_05907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12661__I0 (.I(_05918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12656__I0 (.I(_05918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12651__I0 (.I(_05918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12645__I0 (.I(_05918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12782__I (.I(_05919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12731__I (.I(_05919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12673__I (.I(_05919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12643__I (.I(_05919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12648__S (.I(_05921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12645__S (.I(_05921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12663__I0 (.I(_05923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12658__I0 (.I(_05923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12653__I0 (.I(_05923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12648__I0 (.I(_05923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12698__I0 (.I(_05934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12680__I0 (.I(_05934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12675__I0 (.I(_05934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12667__I0 (.I(_05934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12762__I (.I(_05937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12740__I (.I(_05937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12712__I (.I(_05937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12670__I (.I(_05937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12700__I0 (.I(_05938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12682__I0 (.I(_05938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12677__I0 (.I(_05938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12671__I0 (.I(_05938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12677__S (.I(_05941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12675__S (.I(_05941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12689__S (.I(_05947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12687__A2 (.I(_05947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12686__A2 (.I(_05947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13106__A1 (.I(_05948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13060__A1 (.I(_05948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12807__A1 (.I(_05948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12686__A1 (.I(_05948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12724__I1 (.I(_05950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12705__I1 (.I(_05950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12695__I1 (.I(_05950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12689__I1 (.I(_05950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12770__A2 (.I(_05952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12721__A2 (.I(_05952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12692__A2 (.I(_05952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12695__S (.I(_05953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12693__S (.I(_05953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12705__S (.I(_05959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12703__S (.I(_05959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12733__I0 (.I(_05963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12727__I0 (.I(_05963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12716__I0 (.I(_05963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12710__I0 (.I(_05963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12735__I0 (.I(_05966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12729__I0 (.I(_05966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12718__I0 (.I(_05966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12713__I0 (.I(_05966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13076__I1 (.I(_05971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12916__I1 (.I(_05971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12771__I1 (.I(_05971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12722__I1 (.I(_05971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12757__I0 (.I(_05984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12751__I0 (.I(_05984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12746__I0 (.I(_05984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12741__I0 (.I(_05984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12746__S (.I(_05986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12745__A2 (.I(_05986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12744__A2 (.I(_05986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12751__S (.I(_05989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12750__A2 (.I(_05989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12749__A2 (.I(_05989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12777__I0 (.I(_05992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12766__I0 (.I(_05992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12760__I0 (.I(_05992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12755__I0 (.I(_05992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12757__S (.I(_05993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12755__S (.I(_05993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12763__S (.I(_05996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12760__S (.I(_05996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12786__I0 (.I(_05998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12779__I0 (.I(_05998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12768__I0 (.I(_05998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12763__I0 (.I(_05998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12768__S (.I(_06000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12766__S (.I(_06000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13062__I1 (.I(_06005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12918__I1 (.I(_06005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12809__I1 (.I(_06005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12774__I1 (.I(_06005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12779__S (.I(_06007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12777__S (.I(_06007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12802__I0 (.I(_06010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12797__I0 (.I(_06010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12789__I0 (.I(_06010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12784__I0 (.I(_06010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13412__A2 (.I(_06011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12801__A2 (.I(_06011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12788__A2 (.I(_06011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12783__A2 (.I(_06011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12786__S (.I(_06012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12784__S (.I(_06012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13927__I (.I(_06017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13101__I (.I(_06017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12923__I (.I(_06017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12792__I (.I(_06017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12895__I (.I(_06018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12871__I (.I(_06018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12822__I (.I(_06018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12793__I (.I(_06018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12816__I0 (.I(_06019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12804__I0 (.I(_06019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12799__I0 (.I(_06019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12794__I0 (.I(_06019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12804__S (.I(_06024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12802__S (.I(_06024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12809__S (.I(_06027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12808__A2 (.I(_06027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12807__A2 (.I(_06027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12816__S (.I(_06031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12815__A2 (.I(_06031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12814__A2 (.I(_06031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13088__A1 (.I(_06032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13048__A1 (.I(_06032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12826__A1 (.I(_06032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12814__A1 (.I(_06032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12869__I0 (.I(_06035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12840__I0 (.I(_06035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12831__I0 (.I(_06035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12820__I0 (.I(_06035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12842__I0 (.I(_06038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12833__I0 (.I(_06038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12828__I0 (.I(_06038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12823__I0 (.I(_06038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12828__S (.I(_06040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12827__A2 (.I(_06040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12826__A2 (.I(_06040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14200__A1 (.I(_06046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14166__I (.I(_06046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12866__B (.I(_06046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12836__I (.I(_06046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14206__A1 (.I(_06047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14170__A1 (.I(_06047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13172__A1 (.I(_06047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12837__A1 (.I(_06047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12899__A2 (.I(_06048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12892__A2 (.I(_06048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12881__A2 (.I(_06048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12839__A2 (.I(_06048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12851__A1 (.I(_06052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12848__A1 (.I(_06052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12846__A2 (.I(_06052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12845__A2 (.I(_06052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14201__B (.I(_06056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14157__A1 (.I(_06056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12981__B (.I(_06056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12853__I (.I(_06056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14196__A1 (.I(_06057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14155__A1 (.I(_06057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12937__A1 (.I(_06057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12854__A1 (.I(_06057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14163__A1 (.I(_06062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12991__A1 (.I(_06062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12933__A1 (.I(_06062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12862__I (.I(_06062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14154__I (.I(_06063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12986__A1 (.I(_06063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12936__B2 (.I(_06063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12865__A1 (.I(_06063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13906__A1 (.I(_06065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13784__A1 (.I(_06065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13754__C (.I(_06065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12865__A2 (.I(_06065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12890__I0 (.I(_06070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12884__I0 (.I(_06070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12879__I0 (.I(_06070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12872__I0 (.I(_06070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13024__I (.I(_06072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12927__I (.I(_06072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12898__I (.I(_06072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12875__I (.I(_06072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12893__I0 (.I(_06073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12888__I0 (.I(_06073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12882__I0 (.I(_06073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12877__I0 (.I(_06073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13025__A2 (.I(_06080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13012__A2 (.I(_06080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13007__A2 (.I(_06080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12887__A2 (.I(_06080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12913__I0 (.I(_06086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12908__I0 (.I(_06086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12902__I0 (.I(_06086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12896__I0 (.I(_06086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12921__I0 (.I(_06088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12911__I0 (.I(_06088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12906__I0 (.I(_06088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12900__I0 (.I(_06088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13064__A2 (.I(_06092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13041__A2 (.I(_06092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13030__A2 (.I(_06092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12905__A2 (.I(_06092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13015__I0 (.I(_06105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13010__I0 (.I(_06105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12931__I0 (.I(_06105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12925__I0 (.I(_06105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13019__I0 (.I(_06107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13013__I0 (.I(_06107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13008__I0 (.I(_06107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12929__I0 (.I(_06107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13000__A1 (.I(_06113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12985__A1 (.I(_06113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12936__B1 (.I(_06113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13279__I (.I(_06116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13190__A1 (.I(_06116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12950__A1 (.I(_06116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12940__S (.I(_06116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13209__A1 (.I(_06117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12941__I (.I(_06117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13304__A1 (.I(_06118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13213__I (.I(_06118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13203__A1 (.I(_06118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12944__A1 (.I(_06118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13270__I (.I(_06120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12944__A2 (.I(_06120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13344__I (.I(_06121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12956__A1 (.I(_06121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13290__S (.I(_06122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13220__A1 (.I(_06122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13179__A1 (.I(_06122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12948__A1 (.I(_06122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13942__A1 (.I(_06123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13718__A2 (.I(_06123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13220__A2 (.I(_06123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12948__A2 (.I(_06123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13337__I (.I(_06125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12954__A1 (.I(_06125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12953__A1 (.I(_06125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13261__A1 (.I(_06126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13195__A1 (.I(_06126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13185__S (.I(_06126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12951__A1 (.I(_06126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12954__A2 (.I(_06128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12952__I (.I(_06128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13867__C (.I(_06131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13358__B (.I(_06131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12955__I (.I(_06131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13334__I (.I(_06133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13230__A2 (.I(_06133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12957__A2 (.I(_06133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13664__C (.I(_06134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13311__I (.I(_06134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12958__I (.I(_06134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13902__C2 (.I(_06135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13831__A1 (.I(_06135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13712__C (.I(_06135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12965__A1 (.I(_06135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12960__A3 (.I(_06136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13643__B (.I(_06137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13230__A1 (.I(_06137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12961__I (.I(_06137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13744__A2 (.I(_06139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13380__A1 (.I(_06139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13226__A1 (.I(_06139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12963__I (.I(_06139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13903__A2 (.I(_06140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13899__A2 (.I(_06140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13173__A2 (.I(_06140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12964__A2 (.I(_06140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13506__A1 (.I(_06142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12972__A1 (.I(_06142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12971__A2 (.I(_06142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12968__A1 (.I(_06142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14202__A2 (.I(_06151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14201__A2 (.I(_06151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14200__A2 (.I(_06151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12980__A3 (.I(_06151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14204__A1 (.I(_06153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14159__A1 (.I(_06153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13933__A1 (.I(_06153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12979__A3 (.I(_06153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14168__A2 (.I(_06166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13922__A1 (.I(_06166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13000__A2 (.I(_06166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12997__A1 (.I(_06166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13022__S (.I(_06182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13019__S (.I(_06182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13039__I0 (.I(_06184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13033__I0 (.I(_06184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13028__I0 (.I(_06184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13022__I0 (.I(_06184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13042__I0 (.I(_06186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13037__I0 (.I(_06186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13031__I0 (.I(_06186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13026__I0 (.I(_06186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13235__A2 (.I(_06193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13069__A2 (.I(_06193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13054__A2 (.I(_06193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13036__A2 (.I(_06193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13067__I0 (.I(_06199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13057__I0 (.I(_06199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13050__I0 (.I(_06199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13045__I0 (.I(_06199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13050__S (.I(_06201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13049__A2 (.I(_06201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13048__A2 (.I(_06201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13251__I (.I(_06204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13163__I (.I(_06204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13092__I (.I(_06204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13053__I (.I(_06204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13083__I0 (.I(_06205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13070__I0 (.I(_06205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13065__I0 (.I(_06205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13055__I0 (.I(_06205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13062__S (.I(_06209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13061__A2 (.I(_06209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13060__A2 (.I(_06209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13096__I0 (.I(_06217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13090__I0 (.I(_06217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13085__I0 (.I(_06217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13073__I0 (.I(_06217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13079__S (.I(_06219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13076__S (.I(_06219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14210__I1 (.I(_06221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13603__I1 (.I(_06221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13108__I1 (.I(_06221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13079__I1 (.I(_06221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13892__A2 (.I(_06223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13110__A2 (.I(_06223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13098__A2 (.I(_06223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13082__A2 (.I(_06223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13085__S (.I(_06224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13083__S (.I(_06224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13090__S (.I(_06227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13089__A2 (.I(_06227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13088__A2 (.I(_06227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13116__I0 (.I(_06230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13111__I0 (.I(_06230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13099__I0 (.I(_06230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13094__I0 (.I(_06230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13096__S (.I(_06231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13094__S (.I(_06231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13103__S (.I(_06234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13099__S (.I(_06234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13124__I0 (.I(_06237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13118__I0 (.I(_06237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13113__I0 (.I(_06237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13103__I0 (.I(_06237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13108__S (.I(_06239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13107__A2 (.I(_06239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13106__A2 (.I(_06239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13925__A1 (.I(_06249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13621__A1 (.I(_06249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13616__A1 (.I(_06249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13122__A1 (.I(_06249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13154__I (.I(_06252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13145__I (.I(_06252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13136__I (.I(_06252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13127__I (.I(_06252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13247__I0 (.I(_06273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13242__I0 (.I(_06273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13236__I0 (.I(_06273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13165__I0 (.I(_06273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13249__I0 (.I(_06276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13244__I0 (.I(_06276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13238__I0 (.I(_06276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13168__I0 (.I(_06276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13751__B2 (.I(_06281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13294__A1 (.I(_06281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13188__A3 (.I(_06281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13175__I (.I(_06281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13865__A1 (.I(_06282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13673__B (.I(_06282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13189__A1 (.I(_06282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13176__I (.I(_06282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13869__A4 (.I(_06283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13828__A1 (.I(_06283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13753__B1 (.I(_06283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13200__A1 (.I(_06283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13630__A2 (.I(_06284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13294__A2 (.I(_06284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13187__I (.I(_06284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13178__I (.I(_06284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13886__A2 (.I(_06285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13398__I (.I(_06285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13200__A2 (.I(_06285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13189__C (.I(_06285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13774__A1 (.I(_06289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13648__A1 (.I(_06289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13298__A1 (.I(_06289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13189__A2 (.I(_06289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13856__A2 (.I(_06292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13687__A1 (.I(_06292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13372__I (.I(_06292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13186__I (.I(_06292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13304__A2 (.I(_06300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13276__I (.I(_06300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13209__A2 (.I(_06300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13194__A2 (.I(_06300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13674__A1 (.I(_06304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13655__A1 (.I(_06304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13328__A2 (.I(_06304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13198__A2 (.I(_06304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13696__A2 (.I(_06306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13674__C2 (.I(_06306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13278__A1 (.I(_06306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13200__C (.I(_06306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13773__A1 (.I(_06309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13661__A1 (.I(_06309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13210__A1 (.I(_06309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13203__A2 (.I(_06309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13909__A1 (.I(_06311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13884__A2 (.I(_06311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13820__A1 (.I(_06311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13208__A1 (.I(_06311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13725__B2 (.I(_06314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13720__A2 (.I(_06314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13347__A2 (.I(_06314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13208__A2 (.I(_06314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13352__I (.I(_06316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13330__A1 (.I(_06316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13210__A2 (.I(_06316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13708__A1 (.I(_06318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13333__A1 (.I(_06318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13268__A1 (.I(_06318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13212__I (.I(_06318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13719__I (.I(_06320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13704__C (.I(_06320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13650__A1 (.I(_06320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13214__I (.I(_06320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13796__A1 (.I(_06321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13727__B (.I(_06321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13277__A1 (.I(_06321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13217__A1 (.I(_06321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13827__A2 (.I(_06324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13780__A2 (.I(_06324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13632__A2 (.I(_06324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13218__A4 (.I(_06324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13751__B1 (.I(_06326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13366__A1 (.I(_06326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13332__A2 (.I(_06326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13224__A2 (.I(_06326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13299__I (.I(_06328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13282__A1 (.I(_06328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13222__A1 (.I(_06328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13395__A2 (.I(_06329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13267__I (.I(_06329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13223__I (.I(_06329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13751__C (.I(_06330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13366__B (.I(_06330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13332__B (.I(_06330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13224__B (.I(_06330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13821__B (.I(_06332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13806__B2 (.I(_06332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13629__I (.I(_06332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13226__A2 (.I(_06332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13855__S (.I(_06335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13829__S (.I(_06335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13749__A1 (.I(_06335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13229__S (.I(_06335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13744__B1 (.I(_06338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13665__A1 (.I(_06338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13313__A1 (.I(_06338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13232__I (.I(_06338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13830__C2 (.I(_06339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13799__A1 (.I(_06339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13322__B1 (.I(_06339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13233__B2 (.I(_06339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13238__S (.I(_06341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13236__S (.I(_06341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13418__I0 (.I(_06351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13413__I0 (.I(_06351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13408__I0 (.I(_06351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13253__I0 (.I(_06351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13256__S (.I(_06352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13253__S (.I(_06352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13420__I0 (.I(_06354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13415__I0 (.I(_06354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13410__I0 (.I(_06354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13256__I0 (.I(_06354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13275__A2 (.I(_06360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13263__A2 (.I(_06360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13819__A1 (.I(_06363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13712__A1 (.I(_06363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13710__A2 (.I(_06363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13313__A2 (.I(_06363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13868__I (.I(_06365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13757__C (.I(_06365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13708__C (.I(_06365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13268__B (.I(_06365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13844__A1 (.I(_06367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13684__I (.I(_06367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13285__A1 (.I(_06367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13271__A1 (.I(_06367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13858__A2 (.I(_06370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13674__A2 (.I(_06370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13331__A2 (.I(_06370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13278__B1 (.I(_06370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13703__A1 (.I(_06371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13659__A1 (.I(_06371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13631__A1 (.I(_06371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13274__I (.I(_06371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13820__B2 (.I(_06372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13781__A2 (.I(_06372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13676__B2 (.I(_06372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13278__B2 (.I(_06372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13389__A1 (.I(_06377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13288__A1 (.I(_06377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13287__S (.I(_06377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13280__A1 (.I(_06377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13780__B (.I(_06380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13709__A1 (.I(_06380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13358__A2 (.I(_06380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13283__I (.I(_06380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13781__A1 (.I(_06381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13736__C (.I(_06381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13402__A1 (.I(_06381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13302__B (.I(_06381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13886__A1 (.I(_06382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13724__A1 (.I(_06382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13347__B2 (.I(_06382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13285__A2 (.I(_06382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13912__A3 (.I(_06390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13351__A2 (.I(_06390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13342__A2 (.I(_06390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13298__A2 (.I(_06390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13366__A2 (.I(_06391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13362__I (.I(_06391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13294__A3 (.I(_06391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13797__B2 (.I(_06395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13377__B2 (.I(_06395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13358__A1 (.I(_06395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13298__C (.I(_06395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13856__A1 (.I(_06397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13392__A2 (.I(_06397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13385__A1 (.I(_06397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13300__I (.I(_06397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13913__A1 (.I(_06398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13685__A2 (.I(_06398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13393__A2 (.I(_06398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13301__C (.I(_06398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13313__B1 (.I(_06400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13809__A1 (.I(_06401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13798__A1 (.I(_06401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13348__B2 (.I(_06401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13312__A1 (.I(_06401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13792__B1 (.I(_06402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13661__A3 (.I(_06402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13329__A2 (.I(_06402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13305__I (.I(_06402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13403__A2 (.I(_06403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13373__A2 (.I(_06403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13343__A3 (.I(_06403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13310__A1 (.I(_06403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13778__A1 (.I(_06404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13661__A2 (.I(_06404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13649__I (.I(_06404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13307__A2 (.I(_06404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13794__A2 (.I(_06407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13310__A2 (.I(_06407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13768__B2 (.I(_06411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13317__B1 (.I(_06411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13874__A1 (.I(_06412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13759__C (.I(_06412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13636__I (.I(_06412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13315__I (.I(_06412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13915__A2 (.I(_06413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13405__A2 (.I(_06413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13381__A1 (.I(_06413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13316__A2 (.I(_06413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13771__A1 (.I(_06415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13666__I (.I(_06415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13627__I (.I(_06415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13319__I (.I(_06415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13808__A1 (.I(_06418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13802__A1 (.I(_06418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13343__A2 (.I(_06418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13322__B2 (.I(_06418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13762__B (.I(_06421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13698__A1 (.I(_06421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13678__A1 (.I(_06421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13325__I (.I(_06421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13887__B2 (.I(_06423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13817__A1 (.I(_06423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13742__C (.I(_06423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13336__A1 (.I(_06423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13803__I (.I(_06424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13686__A1 (.I(_06424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13346__I (.I(_06424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13331__A1 (.I(_06424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13792__A1 (.I(_06425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13751__A2 (.I(_06425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13740__A2 (.I(_06425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13329__A1 (.I(_06425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13881__A1 (.I(_06426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13778__B2 (.I(_06426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13356__I (.I(_06426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13330__A2 (.I(_06426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13336__A2 (.I(_06430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13815__I (.I(_06431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13697__A2 (.I(_06431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13675__A1 (.I(_06431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13335__I (.I(_06431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13781__C (.I(_06432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13754__A1 (.I(_06432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13403__A1 (.I(_06432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13336__B (.I(_06432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13662__A1 (.I(_06434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13400__I (.I(_06434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13354__A1 (.I(_06434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13339__A1 (.I(_06434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13846__A1 (.I(_06437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13676__A1 (.I(_06437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13361__A1 (.I(_06437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13343__A1 (.I(_06437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13869__A2 (.I(_06438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13726__A1 (.I(_06438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13401__A1 (.I(_06438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13342__A1 (.I(_06438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13808__B2 (.I(_06442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13736__B2 (.I(_06442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13393__A1 (.I(_06442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13347__A1 (.I(_06442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13909__B1 (.I(_06443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13850__A2 (.I(_06443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13802__B2 (.I(_06443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13347__B1 (.I(_06443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13349__A2 (.I(_06445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13350__C (.I(_06446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13653__A1 (.I(_06447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13386__A2 (.I(_06447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13361__A2 (.I(_06447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13845__B (.I(_06450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13697__B1 (.I(_06450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13355__I (.I(_06450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13918__A1 (.I(_06451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13851__A1 (.I(_06451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13677__A1 (.I(_06451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13357__A2 (.I(_06451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13921__B2 (.I(_06452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13913__A2 (.I(_06452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13805__A2 (.I(_06452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13357__A3 (.I(_06452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13849__B (.I(_06455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13783__B (.I(_06455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13634__I (.I(_06455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13360__I (.I(_06455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13921__A1 (.I(_06456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13743__A2 (.I(_06456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13730__A1 (.I(_06456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13361__C (.I(_06456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13820__A2 (.I(_06458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13740__A3 (.I(_06458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13377__B1 (.I(_06458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13363__I (.I(_06458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13381__A2 (.I(_06461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13902__B2 (.I(_06463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13722__A1 (.I(_06463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13690__A2 (.I(_06463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13371__A1 (.I(_06463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13859__B2 (.I(_06464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13696__B1 (.I(_06464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13377__A2 (.I(_06464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13369__I (.I(_06464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13915__B2 (.I(_06465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13860__A1 (.I(_06465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13819__A2 (.I(_06465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13371__B1 (.I(_06465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13850__A3 (.I(_06466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13820__B1 (.I(_06466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13802__A2 (.I(_06466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13371__B2 (.I(_06466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13921__A2 (.I(_06468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13883__A1 (.I(_06468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13805__A1 (.I(_06468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13373__A1 (.I(_06468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13740__A1 (.I(_06470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13704__A1 (.I(_06470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13392__A1 (.I(_06470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13375__I (.I(_06470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13912__A1 (.I(_06471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13826__A1 (.I(_06471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13713__B1 (.I(_06471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13377__A1 (.I(_06471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13850__A1 (.I(_06472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13753__A2 (.I(_06472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13664__B2 (.I(_06472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13377__C (.I(_06472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13759__B2 (.I(_06475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13721__B (.I(_06475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13683__A2 (.I(_06475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13380__A2 (.I(_06475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13921__C (.I(_06481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13905__A1 (.I(_06481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13397__B1 (.I(_06481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13852__B (.I(_06483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13731__A2 (.I(_06483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13404__A1 (.I(_06483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13396__A1 (.I(_06483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13687__A2 (.I(_06485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13630__A1 (.I(_06485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13394__A1 (.I(_06485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13802__C (.I(_06486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13794__B (.I(_06486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13727__C (.I(_06486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13393__B (.I(_06486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13918__B (.I(_06487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13857__A1 (.I(_06487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13393__C (.I(_06487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13906__A2 (.I(_06490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13826__B (.I(_06490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13675__A2 (.I(_06490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13396__A3 (.I(_06490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13724__A2 (.I(_06493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13707__B1 (.I(_06493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13696__C1 (.I(_06493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13401__A2 (.I(_06493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13780__A1 (.I(_06494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13728__I (.I(_06494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13688__A1 (.I(_06494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13401__B (.I(_06494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13404__A3 (.I(_06497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13406__B1 (.I(_06498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13466__I (.I(_06509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13423__I (.I(_06509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13456__I (.I(_06510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13446__I (.I(_06510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13436__I (.I(_06510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13424__I (.I(_06510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13468__I (.I(_06512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13426__I (.I(_06512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13457__I (.I(_06513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13447__I (.I(_06513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13437__I (.I(_06513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13427__I (.I(_06513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13498__I (.I(_06537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13488__I (.I(_06537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13478__I (.I(_06537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13467__I (.I(_06537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13499__I (.I(_06539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13489__I (.I(_06539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13479__I (.I(_06539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13469__I (.I(_06539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13476__B1 (.I(_06540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13474__B1 (.I(_06540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13472__B1 (.I(_06540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13470__B1 (.I(_06540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13509__A1 (.I(_06562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13507__B (.I(_06562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13511__B2 (.I(_06566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14163__A2 (.I(_06568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13519__A1 (.I(_06568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13515__A2 (.I(_06568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13514__C (.I(_06568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14078__I0 (.I(_06578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14073__I0 (.I(_06578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13893__I0 (.I(_06578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13527__I0 (.I(_06578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13895__I0 (.I(_06581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13623__I0 (.I(_06581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13618__I0 (.I(_06581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13530__I0 (.I(_06581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13560__I (.I(_06583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13551__I (.I(_06583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13542__I (.I(_06583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13533__I (.I(_06583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13540__S (.I(_06584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13538__S (.I(_06584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13536__S (.I(_06584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13534__S (.I(_06584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13576__S (.I(_06604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13574__S (.I(_06604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13572__S (.I(_06604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13570__S (.I(_06604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13603__S (.I(_06621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13601__S (.I(_06621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13917__B (.I(_06640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13888__A2 (.I(_06640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13730__C (.I(_06640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13628__I (.I(_06640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13827__A3 (.I(_06643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13774__B (.I(_06643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13632__A3 (.I(_06643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13705__A2 (.I(_06644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13688__A2 (.I(_06644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13662__A2 (.I(_06644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13632__A4 (.I(_06644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13834__A1 (.I(_06651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13670__A1 (.I(_06651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13700__I (.I(_06655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13646__I (.I(_06655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13644__I (.I(_06655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13756__A2 (.I(_06657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13732__A2 (.I(_06657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13714__A2 (.I(_06657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13670__A2 (.I(_06657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13665__A2 (.I(_06659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13912__A4 (.I(_06660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13905__A2 (.I(_06660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13653__A2 (.I(_06660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13907__A2 (.I(_06661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13674__B2 (.I(_06661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13663__A1 (.I(_06661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13651__A1 (.I(_06661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13846__A2 (.I(_06662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13722__A2 (.I(_06662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13651__A2 (.I(_06662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13777__A1 (.I(_06667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13737__A2 (.I(_06667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13707__A2 (.I(_06667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13658__A1 (.I(_06667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13819__A3 (.I(_06668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13723__A2 (.I(_06668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13657__A2 (.I(_06668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13737__A3 (.I(_06669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13706__I (.I(_06669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13658__A2 (.I(_06669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13885__A2 (.I(_06672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13866__A2 (.I(_06672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13851__A2 (.I(_06672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13664__A1 (.I(_06672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13900__A1 (.I(_06677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13843__A1 (.I(_06677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13668__A1 (.I(_06677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13907__B1 (.I(_06682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13696__B2 (.I(_06682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13686__A2 (.I(_06682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13674__B1 (.I(_06682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13901__B (.I(_06689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13680__A1 (.I(_06689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13902__B1 (.I(_06693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13713__B2 (.I(_06693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13690__A1 (.I(_06693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13869__A1 (.I(_06694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13710__A1 (.I(_06694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13697__A1 (.I(_06694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13685__A1 (.I(_06694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13902__C1 (.I(_06699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13690__B1 (.I(_06699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13890__I (.I(_06704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13862__C (.I(_06704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13713__A2 (.I(_06704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13699__A2 (.I(_06704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13904__A1 (.I(_06707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13699__B (.I(_06707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13759__A2 (.I(_06712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13753__B2 (.I(_06712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13742__A2 (.I(_06712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13712__A2 (.I(_06712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13757__B1 (.I(_06713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13739__A1 (.I(_06713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13725__C (.I(_06713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13708__B1 (.I(_06713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13804__A2 (.I(_06714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13791__A2 (.I(_06714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13776__A2 (.I(_06714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13707__A3 (.I(_06714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13711__A1 (.I(_06716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13730__A2 (.I(_06725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13720__B1 (.I(_06725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13794__A1 (.I(_06726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13753__A1 (.I(_06726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13736__A1 (.I(_06726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13720__A1 (.I(_06726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13885__A1 (.I(_06735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13806__A1 (.I(_06735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13795__B2 (.I(_06735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13729__B2 (.I(_06735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13732__B1 (.I(_06737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13873__A1 (.I(_06739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13849__A1 (.I(_06739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13783__A1 (.I(_06739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13735__A1 (.I(_06739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13744__B2 (.I(_06741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13736__B1 (.I(_06741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13860__A2 (.I(_06744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13778__A2 (.I(_06744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13757__B2 (.I(_06744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13739__A2 (.I(_06744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13822__C (.I(_06753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13785__A2 (.I(_06753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13766__A2 (.I(_06753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13755__A2 (.I(_06753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13755__C (.I(_06759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13759__B1 (.I(_06762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13763__B1 (.I(_06765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13812__A2 (.I(_06772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13800__A2 (.I(_06772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13771__A2 (.I(_06772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13836__A2 (.I(_06774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13801__A2 (.I(_06774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13787__A1 (.I(_06774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13786__A2 (.I(_06774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13820__C (.I(_06776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13805__C (.I(_06776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13793__C (.I(_06776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13775__I (.I(_06776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13819__B (.I(_06779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13805__B1 (.I(_06779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13793__A1 (.I(_06779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13778__B1 (.I(_06779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13784__A2 (.I(_06783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13784__A3 (.I(_06785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13785__B (.I(_06786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13799__A2 (.I(_06790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13797__B1 (.I(_06790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13917__A2 (.I(_06791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13867__B (.I(_06791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13866__A1 (.I(_06791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13791__A1 (.I(_06791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13798__A2 (.I(_06798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13891__B (.I(_06800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13801__B1 (.I(_06800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13801__B2 (.I(_06801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13813__B1 (.I(_06807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13808__B1 (.I(_06807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13814__A1 (.I(_06810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13835__B (.I(_06812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13830__B1 (.I(_06812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13823__B1 (.I(_06812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13813__C1 (.I(_06812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13822__A2 (.I(_06815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13818__A2 (.I(_06816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13822__B2 (.I(_06820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13912__A2 (.I(_06823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13887__A1 (.I(_06823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13867__A1 (.I(_06823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13826__A2 (.I(_06823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13828__A2 (.I(_06824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13834__A2 (.I(_06829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13833__A2 (.I(_06829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13874__A2 (.I(_06834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13841__A2 (.I(_06834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13839__A2 (.I(_06834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13889__A2 (.I(_06836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13863__A2 (.I(_06836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13853__A2 (.I(_06836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13842__A2 (.I(_06836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13876__A2 (.I(_06837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13863__B1 (.I(_06837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13853__B1 (.I(_06837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13842__B1 (.I(_06837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13871__A1 (.I(_06840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13860__B (.I(_06840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13846__B (.I(_06840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13851__B (.I(_06844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13898__B (.I(_06847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13854__A1 (.I(_06847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13862__A2 (.I(_06849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13887__A2 (.I(_06850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13857__A2 (.I(_06850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13861__A1 (.I(_06853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13897__B (.I(_06856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13864__A1 (.I(_06856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13882__A1 (.I(_06858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13866__A3 (.I(_06858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13870__A2 (.I(_06862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13878__B1 (.I(_06866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13886__B1 (.I(_06871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13880__A2 (.I(_06871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13888__B2 (.I(_06879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13901__A2 (.I(_06881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13898__A2 (.I(_06881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13897__A2 (.I(_06881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13891__A2 (.I(_06881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13911__A2 (.I(_06890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13914__A2 (.I(_06892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13923__A2 (.I(_06899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13929__S (.I(_06901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13926__A2 (.I(_06901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13925__A2 (.I(_06901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14086__I0 (.I(_06904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14080__I0 (.I(_06904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14075__I0 (.I(_06904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13929__I0 (.I(_06904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14010__I (.I(_06909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13938__A2 (.I(_06909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13935__I (.I(_06909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13994__I (.I(_06910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13979__I (.I(_06910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13955__I (.I(_06910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13936__I (.I(_06910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14051__I (.I(_06914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14036__I (.I(_06914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13973__I (.I(_06914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13940__B (.I(_06914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14070__B1 (.I(_06919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14065__A2 (.I(_06919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13972__B1 (.I(_06919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13949__B (.I(_06919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13983__A2 (.I(_06938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13980__A2 (.I(_06938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13976__A2 (.I(_06938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13968__A2 (.I(_06938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14069__A2 (.I(_06940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13971__A2 (.I(_06940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14021__I (.I(_06942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14005__I (.I(_06942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13989__I (.I(_06942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13974__I (.I(_06942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13998__A2 (.I(_06952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13995__A2 (.I(_06952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13991__A2 (.I(_06952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13987__A2 (.I(_06952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14048__I (.I(_06963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14033__I (.I(_06963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14018__I (.I(_06963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14002__I (.I(_06963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14015__A2 (.I(_06964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14012__A2 (.I(_06964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14007__A2 (.I(_06964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14003__A2 (.I(_06964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14056__I (.I(_06970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14041__I (.I(_06970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14026__I (.I(_06970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14011__I (.I(_06970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14023__B1 (.I(_06971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14019__B1 (.I(_06971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14015__B1 (.I(_06971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14012__B1 (.I(_06971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14045__A2 (.I(_06987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14042__A2 (.I(_06987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14038__A2 (.I(_06987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14034__A2 (.I(_06987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14047__A2 (.I(_06989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14044__A2 (.I(_06989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14040__A2 (.I(_06989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14037__A2 (.I(_06989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14060__A2 (.I(_06998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14057__A2 (.I(_06998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14053__A2 (.I(_06998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14049__A2 (.I(_06998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14054__A1 (.I(_07001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14070__B2 (.I(_07012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14100__A2 (.I(_07014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14095__A2 (.I(_07014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14083__A2 (.I(_07014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14072__A2 (.I(_07014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14111__I0 (.I(_07021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14101__I0 (.I(_07021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14096__I0 (.I(_07021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14084__I0 (.I(_07021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14183__A1 (.I(_07026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14150__A1 (.I(_07026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14106__A1 (.I(_07026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14090__A1 (.I(_07026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14108__I0 (.I(_07028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14103__I0 (.I(_07028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14098__I0 (.I(_07028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14093__I0 (.I(_07028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14098__S (.I(_07030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14096__S (.I(_07030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14103__S (.I(_07033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14101__S (.I(_07033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14114__S (.I(_07039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14111__S (.I(_07039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14130__I0 (.I(_07041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14125__I0 (.I(_07041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14120__I0 (.I(_07041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14114__I0 (.I(_07041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14133__I0 (.I(_07043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14128__I0 (.I(_07043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14123__I0 (.I(_07043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14118__I0 (.I(_07043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14120__S (.I(_07044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14118__S (.I(_07044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14136__S (.I(_07053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14133__S (.I(_07053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14152__I0 (.I(_07055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14147__I0 (.I(_07055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14142__I0 (.I(_07055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14136__I0 (.I(_07055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14178__I0 (.I(_07057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14172__I0 (.I(_07057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14145__I0 (.I(_07057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14140__I0 (.I(_07057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14167__A2 (.I(_07075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14205__A1 (.I(_07076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14198__A1 (.I(_07076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14195__A1 (.I(_07076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14167__B (.I(_07076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14190__I0 (.I(_07081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14185__I0 (.I(_07081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14180__I0 (.I(_07081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14175__I0 (.I(_07081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14180__S (.I(_07083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14178__S (.I(_07083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14190__S (.I(_07089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14188__S (.I(_07089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14193__A1 (.I(_07092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14220__S (.I(_07106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14218__S (.I(_07106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(io_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(io_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(io_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12934__A3 (.I(\mod.timer_irq ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09111__A2 (.I(\mod.timer_irq ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13558__I0 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13556__I1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09315__A1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13561__I0 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13558__I1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09324__B2 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13570__I0 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13567__I1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09347__B2 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13576__I0 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13574__I1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09362__B2 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13588__I0 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13585__I1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09397__B2 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13590__I0 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13588__I1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09404__A1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13592__I0 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13590__I1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09411__A1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13534__I0 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13520__A1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09244__C2 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13596__A1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13594__I1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09425__A1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13536__I0 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13534__I1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09253__B2 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13998__B2 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13993__A1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09177__I1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14003__B2 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13997__A1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09179__I1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14007__B2 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14000__A1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09181__I1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14015__B2 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14009__A1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09186__I1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09024__I1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14045__B2 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14040__A1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09204__I1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09024__I3 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13965__A1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12458__A1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09156__I (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08978__A2 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13976__B2 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12460__B2 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09159__I1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13983__B2 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13978__A1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09166__I1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09024__I2 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12959__A1 (.I(\mod.u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12448__A1 (.I(\mod.u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09230__I (.I(\mod.u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13174__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09161__I (.I(\mod.u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13995__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13807__I1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13177__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09166__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13998__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13816__I1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13180__A2 (.I(\mod.u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09168__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14003__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13829__I1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13196__A2 (.I(\mod.u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09170__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14015__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13717__A2 (.I(\mod.u_arbiter.i_wb_cpu_rdt[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13128__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09179__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14019__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13734__A2 (.I(\mod.u_arbiter.i_wb_cpu_rdt[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13130__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09181__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14023__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13750__A2 (.I(\mod.u_arbiter.i_wb_cpu_rdt[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13132__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09183__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14027__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13758__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13134__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09186__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13950__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09127__I (.I(\mod.u_arbiter.i_wb_cpu_rdt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14030__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13647__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13137__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09188__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14034__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13848__A2 (.I(\mod.u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13139__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09190__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14038__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13855__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13141__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09192__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14042__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13872__A2 (.I(\mod.u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13143__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09195__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14045__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13879__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13146__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09197__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14049__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13782__A2 (.I(\mod.u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13148__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09199__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14053__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13789__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13150__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09201__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14057__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13807__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13152__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09204__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14060__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13816__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13155__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09206__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14063__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13829__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13157__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09208__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13956__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09132__I (.I(\mod.u_arbiter.i_wb_cpu_rdt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14066__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13229__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13159__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09210__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14069__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13633__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13161__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09213__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13961__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13758__I1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13287__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09137__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13968__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13647__I1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13290__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09143__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13971__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13849__A2 (.I(\mod.u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13183__A2 (.I(\mod.u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09147__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13976__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13855__I1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13185__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09151__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13980__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13873__A2 (.I(\mod.u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13262__A2 (.I(\mod.u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09154__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13983__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13879__I1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13205__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09157__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13987__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13783__A2 (.I(\mod.u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13293__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09159__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09003__I (.I(\mod.u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09000__A2 (.I(\mod.u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08983__A1 (.I(\mod.u_cpu.cpu.branch_op ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08969__A2 (.I(\mod.u_cpu.cpu.branch_op ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07113__I (.I(\mod.u_cpu.cpu.branch_op ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13598__A1 (.I(\mod.u_cpu.cpu.bufreg.i_sh_signed ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13173__A1 (.I(\mod.u_cpu.cpu.bufreg.i_sh_signed ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08996__A2 (.I(\mod.u_cpu.cpu.bufreg.i_sh_signed ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09024__S1 (.I(\mod.u_cpu.cpu.bufreg.lsb[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09011__A1 (.I(\mod.u_cpu.cpu.bufreg.lsb[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08974__I (.I(\mod.u_cpu.cpu.bufreg.lsb[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13933__A2 (.I(\mod.u_cpu.cpu.bufreg.lsb[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13932__A2 (.I(\mod.u_cpu.cpu.bufreg.lsb[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09091__I (.I(\mod.u_cpu.cpu.bufreg.lsb[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09024__S0 (.I(\mod.u_cpu.cpu.bufreg.lsb[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09034__I (.I(\mod.u_cpu.cpu.bufreg2.i_cnt_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08971__A1 (.I(\mod.u_cpu.cpu.bufreg2.i_cnt_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08970__A1 (.I(\mod.u_cpu.cpu.bufreg2.i_cnt_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08982__A2 (.I(\mod.u_cpu.cpu.csr_d_sel ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08969__A3 (.I(\mod.u_cpu.cpu.csr_d_sel ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07121__I (.I(\mod.u_cpu.cpu.csr_d_sel ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07111__A3 (.I(\mod.u_cpu.cpu.csr_d_sel ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09061__I (.I(\mod.u_cpu.cpu.csr_imm ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09057__A2 (.I(\mod.u_cpu.cpu.csr_imm ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07110__A2 (.I(\mod.u_cpu.cpu.csr_imm ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12964__A1 (.I(\mod.u_cpu.cpu.ctrl.i_iscomp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09017__A2 (.I(\mod.u_cpu.cpu.ctrl.i_iscomp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09016__A2 (.I(\mod.u_cpu.cpu.ctrl.i_iscomp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09321__A1 (.I(\mod.u_cpu.cpu.ctrl.o_ibus_adr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09297__A1 (.I(\mod.u_cpu.cpu.ctrl.o_ibus_adr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09295__I (.I(\mod.u_cpu.cpu.ctrl.o_ibus_adr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13448__A1 (.I(\mod.u_cpu.cpu.ctrl.o_ibus_adr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13444__B2 (.I(\mod.u_cpu.cpu.ctrl.o_ibus_adr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09284__A1 (.I(\mod.u_cpu.cpu.ctrl.o_ibus_adr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09279__A1 (.I(\mod.u_cpu.cpu.ctrl.o_ibus_adr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13190__A2 (.I(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13159__I1 (.I(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12940__I1 (.I(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13192__I1 (.I(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13161__I1 (.I(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12942__A2 (.I(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13287__I1 (.I(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13134__I1 (.I(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13184__A2 (.I(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13139__I1 (.I(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08980__A3 (.I(\mod.u_cpu.cpu.genblk3.csr.o_new_irq ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07125__I (.I(\mod.u_cpu.cpu.genblk3.csr.o_new_irq ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10035__A1 (.I(\mod.u_cpu.cpu.immdec.imm11_7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09433__I (.I(\mod.u_cpu.cpu.immdec.imm11_7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10859__A1 (.I(\mod.u_cpu.cpu.immdec.imm11_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09499__A1 (.I(\mod.u_cpu.cpu.immdec.imm11_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09431__I (.I(\mod.u_cpu.cpu.immdec.imm11_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10160__I (.I(\mod.u_cpu.cpu.immdec.imm11_7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09499__A2 (.I(\mod.u_cpu.cpu.immdec.imm11_7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09434__I (.I(\mod.u_cpu.cpu.immdec.imm11_7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13715__I (.I(\mod.u_cpu.cpu.immdec.imm19_12_20[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13713__A1 (.I(\mod.u_cpu.cpu.immdec.imm19_12_20[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07141__A2 (.I(\mod.u_cpu.cpu.immdec.imm19_12_20[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13746__A1 (.I(\mod.u_cpu.cpu.immdec.imm19_12_20[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13731__A1 (.I(\mod.u_cpu.cpu.immdec.imm19_12_20[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07164__A2 (.I(\mod.u_cpu.cpu.immdec.imm19_12_20[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13744__A1 (.I(\mod.u_cpu.cpu.immdec.imm19_12_20[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07171__I (.I(\mod.u_cpu.cpu.immdec.imm19_12_20[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07161__A2 (.I(\mod.u_cpu.cpu.immdec.imm19_12_20[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13764__I0 (.I(\mod.u_cpu.cpu.immdec.imm19_12_20[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13755__A1 (.I(\mod.u_cpu.cpu.immdec.imm19_12_20[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07159__A2 (.I(\mod.u_cpu.cpu.immdec.imm19_12_20[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13842__A1 (.I(\mod.u_cpu.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13762__A2 (.I(\mod.u_cpu.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08968__B (.I(\mod.u_cpu.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07134__A1 (.I(\mod.u_cpu.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13877__A1 (.I(\mod.u_cpu.cpu.immdec.imm24_20[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13863__B2 (.I(\mod.u_cpu.cpu.immdec.imm24_20[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07172__A1 (.I(\mod.u_cpu.cpu.immdec.imm24_20[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07161__B2 (.I(\mod.u_cpu.cpu.immdec.imm24_20[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13760__A1 (.I(\mod.u_cpu.cpu.immdec.imm31 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13637__A1 (.I(\mod.u_cpu.cpu.immdec.imm31 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08970__A2 (.I(\mod.u_cpu.cpu.immdec.imm31 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09436__A1 (.I(\mod.u_cpu.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09096__A1 (.I(\mod.u_cpu.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08979__I (.I(\mod.u_cpu.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08978__B (.I(\mod.u_cpu.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13514__A1 (.I(\mod.u_cpu.cpu.state.o_cnt_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09089__A1 (.I(\mod.u_cpu.cpu.state.o_cnt_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09015__I (.I(\mod.u_cpu.cpu.state.o_cnt_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08985__A1 (.I(\mod.u_cpu.cpu.state.o_cnt_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14157__A2 (.I(\mod.u_cpu.cpu.state.o_cnt_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09089__A4 (.I(\mod.u_cpu.cpu.state.o_cnt_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09016__A1 (.I(\mod.u_cpu.cpu.state.o_cnt_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08985__A4 (.I(\mod.u_cpu.cpu.state.o_cnt_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09088__I (.I(\mod.u_cpu.cpu.state.o_cnt_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09040__A1 (.I(\mod.u_cpu.cpu.state.o_cnt_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08985__A3 (.I(\mod.u_cpu.cpu.state.o_cnt_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07252__I (.I(\mod.u_cpu.raddr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07207__I (.I(\mod.u_cpu.raddr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07198__I (.I(\mod.u_cpu.raddr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07186__I (.I(\mod.u_cpu.raddr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07351__I (.I(\mod.u_cpu.raddr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07182__I (.I(\mod.u_cpu.raddr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13076__I0 (.I(\mod.u_cpu.rf_ram.memory[105][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07988__I1 (.I(\mod.u_cpu.rf_ram.memory[105][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13079__I0 (.I(\mod.u_cpu.rf_ram.memory[105][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08750__I1 (.I(\mod.u_cpu.rf_ram.memory[105][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13042__I1 (.I(\mod.u_cpu.rf_ram.memory[107][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07988__I3 (.I(\mod.u_cpu.rf_ram.memory[107][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13045__I1 (.I(\mod.u_cpu.rf_ram.memory[107][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08750__I3 (.I(\mod.u_cpu.rf_ram.memory[107][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13031__I1 (.I(\mod.u_cpu.rf_ram.memory[108][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07993__A2 (.I(\mod.u_cpu.rf_ram.memory[108][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13033__I1 (.I(\mod.u_cpu.rf_ram.memory[108][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08747__A2 (.I(\mod.u_cpu.rf_ram.memory[108][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12239__I0 (.I(\mod.u_cpu.rf_ram.memory[109][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08746__I (.I(\mod.u_cpu.rf_ram.memory[109][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14101__I1 (.I(\mod.u_cpu.rf_ram.memory[110][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07999__A2 (.I(\mod.u_cpu.rf_ram.memory[110][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14133__I1 (.I(\mod.u_cpu.rf_ram.memory[115][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08016__I3 (.I(\mod.u_cpu.rf_ram.memory[115][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12667__I1 (.I(\mod.u_cpu.rf_ram.memory[121][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08004__I1 (.I(\mod.u_cpu.rf_ram.memory[121][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12671__I1 (.I(\mod.u_cpu.rf_ram.memory[121][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08762__I1 (.I(\mod.u_cpu.rf_ram.memory[121][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12355__I1 (.I(\mod.u_cpu.rf_ram.memory[122][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08004__I2 (.I(\mod.u_cpu.rf_ram.memory[122][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12357__I1 (.I(\mod.u_cpu.rf_ram.memory[122][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08762__I2 (.I(\mod.u_cpu.rf_ram.memory[122][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13530__I1 (.I(\mod.u_cpu.rf_ram.memory[129][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08608__I1 (.I(\mod.u_cpu.rf_ram.memory[129][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12774__I0 (.I(\mod.u_cpu.rf_ram.memory[133][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08612__I1 (.I(\mod.u_cpu.rf_ram.memory[133][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12716__I1 (.I(\mod.u_cpu.rf_ram.memory[138][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07756__I2 (.I(\mod.u_cpu.rf_ram.memory[138][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12718__I1 (.I(\mod.u_cpu.rf_ram.memory[138][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08617__I2 (.I(\mod.u_cpu.rf_ram.memory[138][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12637__I1 (.I(\mod.u_cpu.rf_ram.memory[148][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07752__I0 (.I(\mod.u_cpu.rf_ram.memory[148][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12632__I1 (.I(\mod.u_cpu.rf_ram.memory[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08081__I2 (.I(\mod.u_cpu.rf_ram.memory[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12634__I1 (.I(\mod.u_cpu.rf_ram.memory[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08812__I2 (.I(\mod.u_cpu.rf_ram.memory[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12571__I1 (.I(\mod.u_cpu.rf_ram.memory[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08081__I3 (.I(\mod.u_cpu.rf_ram.memory[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12575__I1 (.I(\mod.u_cpu.rf_ram.memory[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08812__I3 (.I(\mod.u_cpu.rf_ram.memory[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11934__I0 (.I(\mod.u_cpu.rf_ram.memory[169][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07800__I1 (.I(\mod.u_cpu.rf_ram.memory[169][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11936__I0 (.I(\mod.u_cpu.rf_ram.memory[169][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08638__I1 (.I(\mod.u_cpu.rf_ram.memory[169][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12438__I1 (.I(\mod.u_cpu.rf_ram.memory[172][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07806__A2 (.I(\mod.u_cpu.rf_ram.memory[172][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12440__I1 (.I(\mod.u_cpu.rf_ram.memory[172][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08641__A2 (.I(\mod.u_cpu.rf_ram.memory[172][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12435__I0 (.I(\mod.u_cpu.rf_ram.memory[173][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08639__I (.I(\mod.u_cpu.rf_ram.memory[173][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12323__I1 (.I(\mod.u_cpu.rf_ram.memory[179][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07773__I3 (.I(\mod.u_cpu.rf_ram.memory[179][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12375__I1 (.I(\mod.u_cpu.rf_ram.memory[17][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08096__I1 (.I(\mod.u_cpu.rf_ram.memory[17][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12329__I1 (.I(\mod.u_cpu.rf_ram.memory[184][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07786__I0 (.I(\mod.u_cpu.rf_ram.memory[184][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12331__I1 (.I(\mod.u_cpu.rf_ram.memory[184][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08632__I0 (.I(\mod.u_cpu.rf_ram.memory[184][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12318__I1 (.I(\mod.u_cpu.rf_ram.memory[189][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07791__I1 (.I(\mod.u_cpu.rf_ram.memory[189][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12320__I1 (.I(\mod.u_cpu.rf_ram.memory[189][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08634__I1 (.I(\mod.u_cpu.rf_ram.memory[189][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12243__I1 (.I(\mod.u_cpu.rf_ram.memory[196][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07852__A2 (.I(\mod.u_cpu.rf_ram.memory[196][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12245__I1 (.I(\mod.u_cpu.rf_ram.memory[196][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08697__A2 (.I(\mod.u_cpu.rf_ram.memory[196][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12215__I1 (.I(\mod.u_cpu.rf_ram.memory[198][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07857__A2 (.I(\mod.u_cpu.rf_ram.memory[198][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12217__I1 (.I(\mod.u_cpu.rf_ram.memory[198][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08700__A2 (.I(\mod.u_cpu.rf_ram.memory[198][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12198__I0 (.I(\mod.u_cpu.rf_ram.memory[201][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07865__I1 (.I(\mod.u_cpu.rf_ram.memory[201][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12195__I1 (.I(\mod.u_cpu.rf_ram.memory[202][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08691__I2 (.I(\mod.u_cpu.rf_ram.memory[202][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12178__I1 (.I(\mod.u_cpu.rf_ram.memory[204][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07870__A2 (.I(\mod.u_cpu.rf_ram.memory[204][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12180__I1 (.I(\mod.u_cpu.rf_ram.memory[204][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08688__A2 (.I(\mod.u_cpu.rf_ram.memory[204][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12154__I1 (.I(\mod.u_cpu.rf_ram.memory[206][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07875__A2 (.I(\mod.u_cpu.rf_ram.memory[206][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12130__I1 (.I(\mod.u_cpu.rf_ram.memory[208][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07909__A2 (.I(\mod.u_cpu.rf_ram.memory[208][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12132__I1 (.I(\mod.u_cpu.rf_ram.memory[208][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08681__A2 (.I(\mod.u_cpu.rf_ram.memory[208][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12123__I1 (.I(\mod.u_cpu.rf_ram.memory[20][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08101__A2 (.I(\mod.u_cpu.rf_ram.memory[20][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12126__I1 (.I(\mod.u_cpu.rf_ram.memory[20][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08827__A2 (.I(\mod.u_cpu.rf_ram.memory[20][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12117__I1 (.I(\mod.u_cpu.rf_ram.memory[210][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07905__A2 (.I(\mod.u_cpu.rf_ram.memory[210][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12081__I1 (.I(\mod.u_cpu.rf_ram.memory[212][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07919__A2 (.I(\mod.u_cpu.rf_ram.memory[212][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12083__I1 (.I(\mod.u_cpu.rf_ram.memory[212][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08674__A2 (.I(\mod.u_cpu.rf_ram.memory[212][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12018__I1 (.I(\mod.u_cpu.rf_ram.memory[214][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07915__A2 (.I(\mod.u_cpu.rf_ram.memory[214][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12020__I1 (.I(\mod.u_cpu.rf_ram.memory[214][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08677__A2 (.I(\mod.u_cpu.rf_ram.memory[214][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11985__I1 (.I(\mod.u_cpu.rf_ram.memory[216][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08668__A2 (.I(\mod.u_cpu.rf_ram.memory[216][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11954__I1 (.I(\mod.u_cpu.rf_ram.memory[218][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07892__A2 (.I(\mod.u_cpu.rf_ram.memory[218][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11835__I1 (.I(\mod.u_cpu.rf_ram.memory[228][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07928__A2 (.I(\mod.u_cpu.rf_ram.memory[228][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11837__I1 (.I(\mod.u_cpu.rf_ram.memory[228][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08716__A2 (.I(\mod.u_cpu.rf_ram.memory[228][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11817__I1 (.I(\mod.u_cpu.rf_ram.memory[230][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07931__A2 (.I(\mod.u_cpu.rf_ram.memory[230][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11819__I1 (.I(\mod.u_cpu.rf_ram.memory[230][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08719__A2 (.I(\mod.u_cpu.rf_ram.memory[230][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11773__I1 (.I(\mod.u_cpu.rf_ram.memory[236][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07940__A2 (.I(\mod.u_cpu.rf_ram.memory[236][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11777__I1 (.I(\mod.u_cpu.rf_ram.memory[236][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08707__A2 (.I(\mod.u_cpu.rf_ram.memory[236][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11754__I1 (.I(\mod.u_cpu.rf_ram.memory[238][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07945__A2 (.I(\mod.u_cpu.rf_ram.memory[238][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11756__I1 (.I(\mod.u_cpu.rf_ram.memory[238][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08705__I0 (.I(\mod.u_cpu.rf_ram.memory[238][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11717__I1 (.I(\mod.u_cpu.rf_ram.memory[248][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08732__I0 (.I(\mod.u_cpu.rf_ram.memory[248][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11701__I1 (.I(\mod.u_cpu.rf_ram.memory[252][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07963__A2 (.I(\mod.u_cpu.rf_ram.memory[252][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11703__I1 (.I(\mod.u_cpu.rf_ram.memory[252][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08735__A2 (.I(\mod.u_cpu.rf_ram.memory[252][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11696__I1 (.I(\mod.u_cpu.rf_ram.memory[254][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07967__A2 (.I(\mod.u_cpu.rf_ram.memory[254][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11698__I1 (.I(\mod.u_cpu.rf_ram.memory[254][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08738__A2 (.I(\mod.u_cpu.rf_ram.memory[254][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11657__I1 (.I(\mod.u_cpu.rf_ram.memory[258][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08594__I2 (.I(\mod.u_cpu.rf_ram.memory[258][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11637__I1 (.I(\mod.u_cpu.rf_ram.memory[260][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07706__A2 (.I(\mod.u_cpu.rf_ram.memory[260][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11640__I1 (.I(\mod.u_cpu.rf_ram.memory[260][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08597__A2 (.I(\mod.u_cpu.rf_ram.memory[260][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11624__I1 (.I(\mod.u_cpu.rf_ram.memory[262][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07709__A2 (.I(\mod.u_cpu.rf_ram.memory[262][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11626__I1 (.I(\mod.u_cpu.rf_ram.memory[262][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08600__A2 (.I(\mod.u_cpu.rf_ram.memory[262][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11589__I1 (.I(\mod.u_cpu.rf_ram.memory[268][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07717__A2 (.I(\mod.u_cpu.rf_ram.memory[268][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11591__I1 (.I(\mod.u_cpu.rf_ram.memory[268][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08589__A2 (.I(\mod.u_cpu.rf_ram.memory[268][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11577__I1 (.I(\mod.u_cpu.rf_ram.memory[270][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07723__A2 (.I(\mod.u_cpu.rf_ram.memory[270][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11541__I1 (.I(\mod.u_cpu.rf_ram.memory[276][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07676__A2 (.I(\mod.u_cpu.rf_ram.memory[276][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11543__I1 (.I(\mod.u_cpu.rf_ram.memory[276][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08571__A2 (.I(\mod.u_cpu.rf_ram.memory[276][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11529__I1 (.I(\mod.u_cpu.rf_ram.memory[278][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07679__A2 (.I(\mod.u_cpu.rf_ram.memory[278][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11532__I1 (.I(\mod.u_cpu.rf_ram.memory[278][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08574__A2 (.I(\mod.u_cpu.rf_ram.memory[278][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11525__I1 (.I(\mod.u_cpu.rf_ram.memory[27][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08815__I3 (.I(\mod.u_cpu.rf_ram.memory[27][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11493__I1 (.I(\mod.u_cpu.rf_ram.memory[284][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07693__A2 (.I(\mod.u_cpu.rf_ram.memory[284][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11458__I1 (.I(\mod.u_cpu.rf_ram.memory[28][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08089__A2 (.I(\mod.u_cpu.rf_ram.memory[28][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11460__I1 (.I(\mod.u_cpu.rf_ram.memory[28][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08818__A2 (.I(\mod.u_cpu.rf_ram.memory[28][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11440__I1 (.I(\mod.u_cpu.rf_ram.memory[292][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08540__A2 (.I(\mod.u_cpu.rf_ram.memory[292][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11429__I1 (.I(\mod.u_cpu.rf_ram.memory[294][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08543__A2 (.I(\mod.u_cpu.rf_ram.memory[294][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14078__I1 (.I(\mod.u_cpu.rf_ram.memory[299][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07651__I3 (.I(\mod.u_cpu.rf_ram.memory[299][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14080__I1 (.I(\mod.u_cpu.rf_ram.memory[299][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08535__I3 (.I(\mod.u_cpu.rf_ram.memory[299][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11399__I1 (.I(\mod.u_cpu.rf_ram.memory[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08079__I2 (.I(\mod.u_cpu.rf_ram.memory[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11401__I1 (.I(\mod.u_cpu.rf_ram.memory[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08811__I2 (.I(\mod.u_cpu.rf_ram.memory[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11395__I1 (.I(\mod.u_cpu.rf_ram.memory[300][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08532__A2 (.I(\mod.u_cpu.rf_ram.memory[300][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11380__I1 (.I(\mod.u_cpu.rf_ram.memory[302][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07663__A2 (.I(\mod.u_cpu.rf_ram.memory[302][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11343__I1 (.I(\mod.u_cpu.rf_ram.memory[308][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07629__A2 (.I(\mod.u_cpu.rf_ram.memory[308][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11345__I1 (.I(\mod.u_cpu.rf_ram.memory[308][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08560__A2 (.I(\mod.u_cpu.rf_ram.memory[308][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11336__I1 (.I(\mod.u_cpu.rf_ram.memory[30][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08092__A2 (.I(\mod.u_cpu.rf_ram.memory[30][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11340__I1 (.I(\mod.u_cpu.rf_ram.memory[30][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08821__A2 (.I(\mod.u_cpu.rf_ram.memory[30][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11330__I1 (.I(\mod.u_cpu.rf_ram.memory[310][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07633__A2 (.I(\mod.u_cpu.rf_ram.memory[310][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11332__I1 (.I(\mod.u_cpu.rf_ram.memory[310][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08563__A2 (.I(\mod.u_cpu.rf_ram.memory[310][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11317__I1 (.I(\mod.u_cpu.rf_ram.memory[312][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07609__I0 (.I(\mod.u_cpu.rf_ram.memory[312][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11311__I1 (.I(\mod.u_cpu.rf_ram.memory[313][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07609__I1 (.I(\mod.u_cpu.rf_ram.memory[313][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11294__I1 (.I(\mod.u_cpu.rf_ram.memory[316][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07615__A2 (.I(\mod.u_cpu.rf_ram.memory[316][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11296__I1 (.I(\mod.u_cpu.rf_ram.memory[316][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08551__A2 (.I(\mod.u_cpu.rf_ram.memory[316][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11280__I1 (.I(\mod.u_cpu.rf_ram.memory[318][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07620__A2 (.I(\mod.u_cpu.rf_ram.memory[318][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11282__I1 (.I(\mod.u_cpu.rf_ram.memory[318][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08554__A2 (.I(\mod.u_cpu.rf_ram.memory[318][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11241__I1 (.I(\mod.u_cpu.rf_ram.memory[324][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08504__A2 (.I(\mod.u_cpu.rf_ram.memory[324][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11226__I1 (.I(\mod.u_cpu.rf_ram.memory[326][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08507__A2 (.I(\mod.u_cpu.rf_ram.memory[326][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13601__I0 (.I(\mod.u_cpu.rf_ram.memory[329][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07521__I1 (.I(\mod.u_cpu.rf_ram.memory[329][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11190__I1 (.I(\mod.u_cpu.rf_ram.memory[332][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08495__A2 (.I(\mod.u_cpu.rf_ram.memory[332][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11178__I1 (.I(\mod.u_cpu.rf_ram.memory[334][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08498__A2 (.I(\mod.u_cpu.rf_ram.memory[334][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11169__I1 (.I(\mod.u_cpu.rf_ram.memory[335][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07514__I3 (.I(\mod.u_cpu.rf_ram.memory[335][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13418__I1 (.I(\mod.u_cpu.rf_ram.memory[339][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07537__I3 (.I(\mod.u_cpu.rf_ram.memory[339][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13420__I1 (.I(\mod.u_cpu.rf_ram.memory[339][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08518__I3 (.I(\mod.u_cpu.rf_ram.memory[339][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11142__I1 (.I(\mod.u_cpu.rf_ram.memory[340][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08521__A2 (.I(\mod.u_cpu.rf_ram.memory[340][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11131__I1 (.I(\mod.u_cpu.rf_ram.memory[342][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08524__A2 (.I(\mod.u_cpu.rf_ram.memory[342][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11092__I1 (.I(\mod.u_cpu.rf_ram.memory[348][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08513__A2 (.I(\mod.u_cpu.rf_ram.memory[348][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13165__I1 (.I(\mod.u_cpu.rf_ram.memory[349][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07516__I1 (.I(\mod.u_cpu.rf_ram.memory[349][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11036__I1 (.I(\mod.u_cpu.rf_ram.memory[356][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07597__A2 (.I(\mod.u_cpu.rf_ram.memory[356][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11039__I1 (.I(\mod.u_cpu.rf_ram.memory[356][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08484__A2 (.I(\mod.u_cpu.rf_ram.memory[356][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11022__I1 (.I(\mod.u_cpu.rf_ram.memory[358][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07600__A2 (.I(\mod.u_cpu.rf_ram.memory[358][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11024__I1 (.I(\mod.u_cpu.rf_ram.memory[358][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08487__A2 (.I(\mod.u_cpu.rf_ram.memory[358][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11016__I1 (.I(\mod.u_cpu.rf_ram.memory[35][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08118__I3 (.I(\mod.u_cpu.rf_ram.memory[35][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11018__I1 (.I(\mod.u_cpu.rf_ram.memory[35][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08847__I3 (.I(\mod.u_cpu.rf_ram.memory[35][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11010__I1 (.I(\mod.u_cpu.rf_ram.memory[360][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07584__I0 (.I(\mod.u_cpu.rf_ram.memory[360][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10982__I1 (.I(\mod.u_cpu.rf_ram.memory[364][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07588__A2 (.I(\mod.u_cpu.rf_ram.memory[364][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10969__I1 (.I(\mod.u_cpu.rf_ram.memory[366][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07591__A2 (.I(\mod.u_cpu.rf_ram.memory[366][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10971__I1 (.I(\mod.u_cpu.rf_ram.memory[366][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08478__A2 (.I(\mod.u_cpu.rf_ram.memory[366][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12929__I1 (.I(\mod.u_cpu.rf_ram.memory[369][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07565__I1 (.I(\mod.u_cpu.rf_ram.memory[369][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10950__I1 (.I(\mod.u_cpu.rf_ram.memory[36][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08121__A2 (.I(\mod.u_cpu.rf_ram.memory[36][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10952__I1 (.I(\mod.u_cpu.rf_ram.memory[36][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08850__A2 (.I(\mod.u_cpu.rf_ram.memory[36][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10931__I1 (.I(\mod.u_cpu.rf_ram.memory[372][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07570__A2 (.I(\mod.u_cpu.rf_ram.memory[372][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10933__I1 (.I(\mod.u_cpu.rf_ram.memory[372][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08464__A2 (.I(\mod.u_cpu.rf_ram.memory[372][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10919__I1 (.I(\mod.u_cpu.rf_ram.memory[374][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07575__A2 (.I(\mod.u_cpu.rf_ram.memory[374][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12925__I1 (.I(\mod.u_cpu.rf_ram.memory[379][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08459__I3 (.I(\mod.u_cpu.rf_ram.memory[379][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10886__I1 (.I(\mod.u_cpu.rf_ram.memory[380][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08455__A2 (.I(\mod.u_cpu.rf_ram.memory[380][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10871__I1 (.I(\mod.u_cpu.rf_ram.memory[382][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07560__A2 (.I(\mod.u_cpu.rf_ram.memory[382][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10829__I1 (.I(\mod.u_cpu.rf_ram.memory[388][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07366__I0 (.I(\mod.u_cpu.rf_ram.memory[388][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10832__I1 (.I(\mod.u_cpu.rf_ram.memory[388][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08438__I0 (.I(\mod.u_cpu.rf_ram.memory[388][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10823__I1 (.I(\mod.u_cpu.rf_ram.memory[38][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08124__A2 (.I(\mod.u_cpu.rf_ram.memory[38][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10825__I1 (.I(\mod.u_cpu.rf_ram.memory[38][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08853__A2 (.I(\mod.u_cpu.rf_ram.memory[38][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10818__I1 (.I(\mod.u_cpu.rf_ram.memory[390][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07366__I2 (.I(\mod.u_cpu.rf_ram.memory[390][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10792__I1 (.I(\mod.u_cpu.rf_ram.memory[394][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07376__I2 (.I(\mod.u_cpu.rf_ram.memory[394][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10767__I1 (.I(\mod.u_cpu.rf_ram.memory[398][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07382__I2 (.I(\mod.u_cpu.rf_ram.memory[398][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10761__I1 (.I(\mod.u_cpu.rf_ram.memory[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08079__I3 (.I(\mod.u_cpu.rf_ram.memory[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10763__I1 (.I(\mod.u_cpu.rf_ram.memory[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08811__I3 (.I(\mod.u_cpu.rf_ram.memory[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10756__I1 (.I(\mod.u_cpu.rf_ram.memory[400][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07416__I0 (.I(\mod.u_cpu.rf_ram.memory[400][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10751__I1 (.I(\mod.u_cpu.rf_ram.memory[401][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07416__I1 (.I(\mod.u_cpu.rf_ram.memory[401][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10733__I1 (.I(\mod.u_cpu.rf_ram.memory[404][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08429__A2 (.I(\mod.u_cpu.rf_ram.memory[404][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10719__I1 (.I(\mod.u_cpu.rf_ram.memory[406][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07425__A2 (.I(\mod.u_cpu.rf_ram.memory[406][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10722__I1 (.I(\mod.u_cpu.rf_ram.memory[406][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08432__A2 (.I(\mod.u_cpu.rf_ram.memory[406][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10709__I1 (.I(\mod.u_cpu.rf_ram.memory[408][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07391__I0 (.I(\mod.u_cpu.rf_ram.memory[408][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10711__I1 (.I(\mod.u_cpu.rf_ram.memory[408][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08416__I0 (.I(\mod.u_cpu.rf_ram.memory[408][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10673__I1 (.I(\mod.u_cpu.rf_ram.memory[414][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07407__A2 (.I(\mod.u_cpu.rf_ram.memory[414][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10650__I1 (.I(\mod.u_cpu.rf_ram.memory[418][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08384__I2 (.I(\mod.u_cpu.rf_ram.memory[418][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10636__I1 (.I(\mod.u_cpu.rf_ram.memory[420][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07448__A2 (.I(\mod.u_cpu.rf_ram.memory[420][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10638__I1 (.I(\mod.u_cpu.rf_ram.memory[420][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08388__A2 (.I(\mod.u_cpu.rf_ram.memory[420][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10626__I1 (.I(\mod.u_cpu.rf_ram.memory[422][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07456__A2 (.I(\mod.u_cpu.rf_ram.memory[422][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10628__I1 (.I(\mod.u_cpu.rf_ram.memory[422][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08391__A2 (.I(\mod.u_cpu.rf_ram.memory[422][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10585__I1 (.I(\mod.u_cpu.rf_ram.memory[428][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07469__A2 (.I(\mod.u_cpu.rf_ram.memory[428][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10587__I1 (.I(\mod.u_cpu.rf_ram.memory[428][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08377__A2 (.I(\mod.u_cpu.rf_ram.memory[428][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10582__I1 (.I(\mod.u_cpu.rf_ram.memory[42][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08845__I2 (.I(\mod.u_cpu.rf_ram.memory[42][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10573__I1 (.I(\mod.u_cpu.rf_ram.memory[430][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07476__A2 (.I(\mod.u_cpu.rf_ram.memory[430][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10536__I1 (.I(\mod.u_cpu.rf_ram.memory[436][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07487__A2 (.I(\mod.u_cpu.rf_ram.memory[436][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10538__I1 (.I(\mod.u_cpu.rf_ram.memory[436][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08398__A2 (.I(\mod.u_cpu.rf_ram.memory[436][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10525__I1 (.I(\mod.u_cpu.rf_ram.memory[438][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07490__A2 (.I(\mod.u_cpu.rf_ram.memory[438][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10527__I1 (.I(\mod.u_cpu.rf_ram.memory[438][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08401__A2 (.I(\mod.u_cpu.rf_ram.memory[438][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10517__I1 (.I(\mod.u_cpu.rf_ram.memory[440][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08405__I0 (.I(\mod.u_cpu.rf_ram.memory[440][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10491__I1 (.I(\mod.u_cpu.rf_ram.memory[444][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07497__A2 (.I(\mod.u_cpu.rf_ram.memory[444][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10493__I1 (.I(\mod.u_cpu.rf_ram.memory[444][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08408__A2 (.I(\mod.u_cpu.rf_ram.memory[444][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10477__I1 (.I(\mod.u_cpu.rf_ram.memory[446][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07502__A2 (.I(\mod.u_cpu.rf_ram.memory[446][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10479__I1 (.I(\mod.u_cpu.rf_ram.memory[446][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08411__A2 (.I(\mod.u_cpu.rf_ram.memory[446][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10454__I1 (.I(\mod.u_cpu.rf_ram.memory[44][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08130__A2 (.I(\mod.u_cpu.rf_ram.memory[44][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10458__I1 (.I(\mod.u_cpu.rf_ram.memory[44][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08842__A2 (.I(\mod.u_cpu.rf_ram.memory[44][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10449__I1 (.I(\mod.u_cpu.rf_ram.memory[450][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07194__I2 (.I(\mod.u_cpu.rf_ram.memory[450][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10451__I1 (.I(\mod.u_cpu.rf_ram.memory[450][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08291__I2 (.I(\mod.u_cpu.rf_ram.memory[450][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10443__I1 (.I(\mod.u_cpu.rf_ram.memory[451][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07194__I3 (.I(\mod.u_cpu.rf_ram.memory[451][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10445__I1 (.I(\mod.u_cpu.rf_ram.memory[451][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08291__I3 (.I(\mod.u_cpu.rf_ram.memory[451][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10438__I1 (.I(\mod.u_cpu.rf_ram.memory[452][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07206__A2 (.I(\mod.u_cpu.rf_ram.memory[452][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10440__I1 (.I(\mod.u_cpu.rf_ram.memory[452][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08294__A2 (.I(\mod.u_cpu.rf_ram.memory[452][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10425__I1 (.I(\mod.u_cpu.rf_ram.memory[454][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07218__A2 (.I(\mod.u_cpu.rf_ram.memory[454][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10428__I1 (.I(\mod.u_cpu.rf_ram.memory[454][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08297__A2 (.I(\mod.u_cpu.rf_ram.memory[454][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10414__I1 (.I(\mod.u_cpu.rf_ram.memory[456][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07233__I0 (.I(\mod.u_cpu.rf_ram.memory[456][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10416__I1 (.I(\mod.u_cpu.rf_ram.memory[456][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08288__I0 (.I(\mod.u_cpu.rf_ram.memory[456][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10402__I1 (.I(\mod.u_cpu.rf_ram.memory[458][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07233__I2 (.I(\mod.u_cpu.rf_ram.memory[458][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10404__I1 (.I(\mod.u_cpu.rf_ram.memory[458][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08288__I2 (.I(\mod.u_cpu.rf_ram.memory[458][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10390__I1 (.I(\mod.u_cpu.rf_ram.memory[460][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07236__A2 (.I(\mod.u_cpu.rf_ram.memory[460][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10393__I1 (.I(\mod.u_cpu.rf_ram.memory[460][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08281__A2 (.I(\mod.u_cpu.rf_ram.memory[460][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10375__I1 (.I(\mod.u_cpu.rf_ram.memory[462][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07240__A2 (.I(\mod.u_cpu.rf_ram.memory[462][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10377__I1 (.I(\mod.u_cpu.rf_ram.memory[462][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08279__I0 (.I(\mod.u_cpu.rf_ram.memory[462][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10338__I1 (.I(\mod.u_cpu.rf_ram.memory[468][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07268__A2 (.I(\mod.u_cpu.rf_ram.memory[468][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10340__I1 (.I(\mod.u_cpu.rf_ram.memory[468][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08316__A2 (.I(\mod.u_cpu.rf_ram.memory[468][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10329__I1 (.I(\mod.u_cpu.rf_ram.memory[46][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08133__A2 (.I(\mod.u_cpu.rf_ram.memory[46][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10324__I1 (.I(\mod.u_cpu.rf_ram.memory[470][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07275__A2 (.I(\mod.u_cpu.rf_ram.memory[470][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10326__I1 (.I(\mod.u_cpu.rf_ram.memory[470][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08319__A2 (.I(\mod.u_cpu.rf_ram.memory[470][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10289__I1 (.I(\mod.u_cpu.rf_ram.memory[476][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07251__A2 (.I(\mod.u_cpu.rf_ram.memory[476][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10291__I1 (.I(\mod.u_cpu.rf_ram.memory[476][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08307__A2 (.I(\mod.u_cpu.rf_ram.memory[476][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10273__I1 (.I(\mod.u_cpu.rf_ram.memory[478][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07256__A2 (.I(\mod.u_cpu.rf_ram.memory[478][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10275__I1 (.I(\mod.u_cpu.rf_ram.memory[478][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08310__A2 (.I(\mod.u_cpu.rf_ram.memory[478][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10230__I1 (.I(\mod.u_cpu.rf_ram.memory[484][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07316__A2 (.I(\mod.u_cpu.rf_ram.memory[484][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10232__I1 (.I(\mod.u_cpu.rf_ram.memory[484][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08364__A2 (.I(\mod.u_cpu.rf_ram.memory[484][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10221__I1 (.I(\mod.u_cpu.rf_ram.memory[486][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08368__A2 (.I(\mod.u_cpu.rf_ram.memory[486][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12419__I0 (.I(\mod.u_cpu.rf_ram.memory[489][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08355__I1 (.I(\mod.u_cpu.rf_ram.memory[489][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10199__I1 (.I(\mod.u_cpu.rf_ram.memory[48][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08114__I0 (.I(\mod.u_cpu.rf_ram.memory[48][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10201__I1 (.I(\mod.u_cpu.rf_ram.memory[48][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08836__I0 (.I(\mod.u_cpu.rf_ram.memory[48][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10188__I1 (.I(\mod.u_cpu.rf_ram.memory[490][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07331__I2 (.I(\mod.u_cpu.rf_ram.memory[490][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10182__I1 (.I(\mod.u_cpu.rf_ram.memory[491][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07331__I3 (.I(\mod.u_cpu.rf_ram.memory[491][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10176__I1 (.I(\mod.u_cpu.rf_ram.memory[492][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07334__A2 (.I(\mod.u_cpu.rf_ram.memory[492][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10156__I1 (.I(\mod.u_cpu.rf_ram.memory[494][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07342__A2 (.I(\mod.u_cpu.rf_ram.memory[494][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12370__I1 (.I(\mod.u_cpu.rf_ram.memory[499][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07285__I3 (.I(\mod.u_cpu.rf_ram.memory[499][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12372__I1 (.I(\mod.u_cpu.rf_ram.memory[499][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08327__I3 (.I(\mod.u_cpu.rf_ram.memory[499][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11811__I1 (.I(\mod.u_cpu.rf_ram.memory[49][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08114__I1 (.I(\mod.u_cpu.rf_ram.memory[49][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11813__I1 (.I(\mod.u_cpu.rf_ram.memory[49][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08836__I1 (.I(\mod.u_cpu.rf_ram.memory[49][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10115__I1 (.I(\mod.u_cpu.rf_ram.memory[500][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07288__A2 (.I(\mod.u_cpu.rf_ram.memory[500][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10117__I1 (.I(\mod.u_cpu.rf_ram.memory[500][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08330__A2 (.I(\mod.u_cpu.rf_ram.memory[500][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10102__I1 (.I(\mod.u_cpu.rf_ram.memory[502][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07291__A2 (.I(\mod.u_cpu.rf_ram.memory[502][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10104__I1 (.I(\mod.u_cpu.rf_ram.memory[502][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08334__A2 (.I(\mod.u_cpu.rf_ram.memory[502][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10066__I1 (.I(\mod.u_cpu.rf_ram.memory[507][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07298__I3 (.I(\mod.u_cpu.rf_ram.memory[507][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10061__I1 (.I(\mod.u_cpu.rf_ram.memory[508][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07303__A2 (.I(\mod.u_cpu.rf_ram.memory[508][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10049__I1 (.I(\mod.u_cpu.rf_ram.memory[510][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07308__A2 (.I(\mod.u_cpu.rf_ram.memory[510][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10030__I1 (.I(\mod.u_cpu.rf_ram.memory[512][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08216__I0 (.I(\mod.u_cpu.rf_ram.memory[512][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10014__I1 (.I(\mod.u_cpu.rf_ram.memory[515][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08216__I3 (.I(\mod.u_cpu.rf_ram.memory[515][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09992__I1 (.I(\mod.u_cpu.rf_ram.memory[518][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08230__A2 (.I(\mod.u_cpu.rf_ram.memory[518][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09987__I1 (.I(\mod.u_cpu.rf_ram.memory[51][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08114__I3 (.I(\mod.u_cpu.rf_ram.memory[51][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09989__I1 (.I(\mod.u_cpu.rf_ram.memory[51][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08836__I3 (.I(\mod.u_cpu.rf_ram.memory[51][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09973__I1 (.I(\mod.u_cpu.rf_ram.memory[522][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08909__I2 (.I(\mod.u_cpu.rf_ram.memory[522][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09926__I1 (.I(\mod.u_cpu.rf_ram.memory[52][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08112__I0 (.I(\mod.u_cpu.rf_ram.memory[52][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09928__I1 (.I(\mod.u_cpu.rf_ram.memory[52][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08835__I0 (.I(\mod.u_cpu.rf_ram.memory[52][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09908__I1 (.I(\mod.u_cpu.rf_ram.memory[532][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08257__A2 (.I(\mod.u_cpu.rf_ram.memory[532][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09896__I1 (.I(\mod.u_cpu.rf_ram.memory[534][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08261__A2 (.I(\mod.u_cpu.rf_ram.memory[534][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09862__I1 (.I(\mod.u_cpu.rf_ram.memory[53][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08112__I1 (.I(\mod.u_cpu.rf_ram.memory[53][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09866__I1 (.I(\mod.u_cpu.rf_ram.memory[53][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08835__I1 (.I(\mod.u_cpu.rf_ram.memory[53][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09857__I1 (.I(\mod.u_cpu.rf_ram.memory[540][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08922__A2 (.I(\mod.u_cpu.rf_ram.memory[540][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09847__I1 (.I(\mod.u_cpu.rf_ram.memory[542][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08925__A2 (.I(\mod.u_cpu.rf_ram.memory[542][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09791__I1 (.I(\mod.u_cpu.rf_ram.memory[548][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08152__A2 (.I(\mod.u_cpu.rf_ram.memory[548][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09794__I1 (.I(\mod.u_cpu.rf_ram.memory[548][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08864__A2 (.I(\mod.u_cpu.rf_ram.memory[548][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09727__I1 (.I(\mod.u_cpu.rf_ram.memory[555][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08166__I3 (.I(\mod.u_cpu.rf_ram.memory[555][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09721__I1 (.I(\mod.u_cpu.rf_ram.memory[556][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08873__A2 (.I(\mod.u_cpu.rf_ram.memory[556][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09700__I1 (.I(\mod.u_cpu.rf_ram.memory[558][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08876__A2 (.I(\mod.u_cpu.rf_ram.memory[558][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09689__I1 (.I(\mod.u_cpu.rf_ram.memory[55][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08835__I3 (.I(\mod.u_cpu.rf_ram.memory[55][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09641__I1 (.I(\mod.u_cpu.rf_ram.memory[564][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08204__A2 (.I(\mod.u_cpu.rf_ram.memory[564][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09643__I1 (.I(\mod.u_cpu.rf_ram.memory[564][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08892__A2 (.I(\mod.u_cpu.rf_ram.memory[564][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09623__I1 (.I(\mod.u_cpu.rf_ram.memory[566][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08208__A2 (.I(\mod.u_cpu.rf_ram.memory[566][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09564__I1 (.I(\mod.u_cpu.rf_ram.memory[572][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08191__A2 (.I(\mod.u_cpu.rf_ram.memory[572][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09536__I1 (.I(\mod.u_cpu.rf_ram.memory[574][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08195__A2 (.I(\mod.u_cpu.rf_ram.memory[574][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09542__I1 (.I(\mod.u_cpu.rf_ram.memory[574][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08886__A2 (.I(\mod.u_cpu.rf_ram.memory[574][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12111__I1 (.I(\mod.u_cpu.rf_ram.memory[68][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08047__A2 (.I(\mod.u_cpu.rf_ram.memory[68][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12113__I1 (.I(\mod.u_cpu.rf_ram.memory[68][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08801__A2 (.I(\mod.u_cpu.rf_ram.memory[68][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11854__I1 (.I(\mod.u_cpu.rf_ram.memory[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08076__I2 (.I(\mod.u_cpu.rf_ram.memory[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11857__I1 (.I(\mod.u_cpu.rf_ram.memory[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08810__I2 (.I(\mod.u_cpu.rf_ram.memory[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11864__I1 (.I(\mod.u_cpu.rf_ram.memory[70][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08052__A2 (.I(\mod.u_cpu.rf_ram.memory[70][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11866__I1 (.I(\mod.u_cpu.rf_ram.memory[70][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08804__A2 (.I(\mod.u_cpu.rf_ram.memory[70][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11871__I1 (.I(\mod.u_cpu.rf_ram.memory[72][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08796__I0 (.I(\mod.u_cpu.rf_ram.memory[72][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12173__I1 (.I(\mod.u_cpu.rf_ram.memory[76][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08064__A2 (.I(\mod.u_cpu.rf_ram.memory[76][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12175__I1 (.I(\mod.u_cpu.rf_ram.memory[76][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08793__A2 (.I(\mod.u_cpu.rf_ram.memory[76][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12710__I1 (.I(\mod.u_cpu.rf_ram.memory[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08076__I3 (.I(\mod.u_cpu.rf_ram.memory[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14114__I1 (.I(\mod.u_cpu.rf_ram.memory[87][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08784__I3 (.I(\mod.u_cpu.rf_ram.memory[87][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14175__I1 (.I(\mod.u_cpu.rf_ram.memory[88][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08786__I0 (.I(\mod.u_cpu.rf_ram.memory[88][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09504__I0 (.I(\mod.u_cpu.rf_ram.memory[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08082__I1 (.I(\mod.u_cpu.rf_ram.memory[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12860__A2 (.I(\mod.u_cpu.rf_ram_if.rtrig1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12859__A1 (.I(\mod.u_cpu.rf_ram_if.rtrig1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08997__S (.I(\mod.u_cpu.rf_ram_if.rtrig1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15315__D (.I(\mod.u_cpu.rf_ram_if.wdata1_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09506__A2 (.I(\mod.u_cpu.rf_ram_if.wdata1_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09317__A2 (.I(\mod.u_scanchain_local.module_data_in[50] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15313__D (.I(\mod.u_scanchain_local.module_data_in[69] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09082__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09105__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09083__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15646__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15645__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15644__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15643__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15642__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15641__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15640__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15639__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15638__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15637__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15636__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15635__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15634__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15633__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15632__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15631__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15630__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15629__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15628__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15627__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15626__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15625__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15624__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15623__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15622__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15621__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15620__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15619__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15618__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15617__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15616__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15615__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15614__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15613__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15612__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15611__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15610__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15609__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15608__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15607__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15606__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15605__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15604__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15603__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15602__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15601__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15600__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15599__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15598__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15597__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15596__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15595__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15594__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15593__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15592__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15591__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15590__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15589__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15588__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15587__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15586__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15585__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15584__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15583__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15582__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15581__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15580__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15579__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15578__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15577__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15576__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15575__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15574__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15573__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15572__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15571__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15570__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15569__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15568__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15567__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15566__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15565__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15564__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15563__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15562__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15561__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15560__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15559__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15558__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15557__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15556__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15555__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15554__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15553__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15552__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15551__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15550__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15549__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15548__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15547__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15546__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15545__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15544__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15543__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15542__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15541__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15540__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15539__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15538__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15537__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15536__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15535__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15534__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15533__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15532__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15531__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15530__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15529__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15528__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15527__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15526__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15525__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15524__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15523__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15522__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15521__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15520__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15519__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15518__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15517__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15516__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15515__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15514__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15513__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15512__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15511__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15510__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15509__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15508__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15507__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15506__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15505__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15504__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15503__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15502__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15501__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15500__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15499__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15498__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15497__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15496__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15495__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15494__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15493__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15492__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15491__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15490__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15489__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15488__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15487__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15486__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15485__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15484__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15483__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15482__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15481__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15480__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15479__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15478__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15477__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15476__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15475__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15474__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15473__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15472__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15471__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15470__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15469__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15468__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15467__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15466__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15465__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15464__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15463__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15462__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15461__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15460__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15459__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15458__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15457__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15456__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15455__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15454__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15453__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15452__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15451__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15450__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15449__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15448__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15447__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15446__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15445__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15444__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15443__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15442__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15441__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15440__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15439__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15438__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15437__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15436__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15435__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15434__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15433__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15432__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15431__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15430__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15429__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15428__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15427__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15426__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15425__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15424__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15423__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15422__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15421__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15420__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15419__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15418__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15417__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15416__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15415__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15414__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15413__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15412__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15411__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15410__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15409__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15408__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15407__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15406__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15405__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15404__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15403__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15402__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15401__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15400__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15399__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15398__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15397__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15396__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15395__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15394__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15393__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15392__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15391__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15390__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15389__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15388__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15387__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15386__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15385__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15384__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15383__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15382__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15381__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15380__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15379__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15378__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15377__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15376__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15375__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15374__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15373__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15372__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15371__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15370__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15369__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15368__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15367__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15366__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15365__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15364__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15363__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15362__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15361__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15360__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15359__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15358__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15357__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15356__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15355__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15354__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15353__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15352__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15351__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15350__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15349__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15348__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15347__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15346__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15345__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15344__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15343__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15342__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15341__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15340__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15339__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15338__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15337__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15336__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15335__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15334__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15333__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15332__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15331__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15330__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15329__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15328__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15327__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15326__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15325__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15324__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15323__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15322__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15321__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15320__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15319__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15318__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15317__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15316__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15315__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15314__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15242__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15241__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15240__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15239__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15238__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15237__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15236__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15235__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15234__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15233__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15232__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15231__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15230__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15229__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15228__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15227__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15226__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15225__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15224__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15223__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15222__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15221__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15220__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15219__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15218__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15217__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15216__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15215__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15214__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15213__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15212__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15211__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15210__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15209__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15208__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15207__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15206__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15205__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15204__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15203__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15202__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15201__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15200__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15199__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15198__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15197__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15196__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15195__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15194__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15193__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15192__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15191__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15190__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15189__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15188__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15187__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15186__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15185__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15184__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15183__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15182__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15181__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15180__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15179__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15178__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15177__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15176__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15175__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15174__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15173__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15172__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15171__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15170__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15169__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15168__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15167__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15166__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15165__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15164__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15163__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15162__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15161__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15160__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15159__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15158__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15157__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15156__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15155__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15154__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15153__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15152__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15151__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15150__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15149__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15148__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15147__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15146__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15145__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15144__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15143__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15142__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15141__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15140__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15139__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15138__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15137__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15136__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15135__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15134__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15133__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15132__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15131__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15130__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15129__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15128__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15127__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15126__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15125__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15124__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15123__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15122__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15121__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15120__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15119__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15118__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15117__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15116__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15115__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15114__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15113__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15112__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15111__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15110__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15109__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15108__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15107__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15106__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15105__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15104__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15103__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15102__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15101__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15100__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15099__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15098__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15097__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15096__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15095__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15094__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15093__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15092__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15091__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15090__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15089__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15088__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15087__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15086__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15085__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15084__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15083__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15082__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15081__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15080__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15079__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15078__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15077__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15076__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15075__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15074__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15073__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15072__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15071__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15070__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15069__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15068__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15067__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15066__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15065__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15064__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15063__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15062__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15061__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15060__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15059__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15058__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15057__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15056__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15055__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15054__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15053__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15052__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15051__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15050__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15049__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15048__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15047__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15046__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15045__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15044__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15043__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15042__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15041__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15040__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15039__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15038__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15037__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15036__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15035__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15034__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15033__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15032__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15031__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15030__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15029__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15028__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15027__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15026__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15025__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15024__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15023__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15022__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15021__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15020__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15019__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15018__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15017__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15016__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15015__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15014__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15013__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15012__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15011__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15010__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15009__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15008__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15007__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15006__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15005__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15004__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15003__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15002__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15001__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15000__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14999__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14998__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14997__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14996__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14995__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14994__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14993__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14992__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14991__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14990__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14989__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14988__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14987__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14986__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14985__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14984__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14983__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14982__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14981__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14980__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14979__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14978__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14977__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14976__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14975__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14974__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14973__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14972__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14971__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14970__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14969__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14968__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14967__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14966__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14965__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14964__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14963__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14962__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14961__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14960__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14959__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14958__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14957__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14956__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14955__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14954__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14953__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14952__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14951__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14950__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14949__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14948__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14947__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14946__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14945__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14944__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14943__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14942__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14941__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14940__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14939__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14938__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14937__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14936__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14935__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14934__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14933__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14932__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14931__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14930__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14929__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14928__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14927__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14926__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14925__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14924__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14923__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14922__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14921__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14920__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14919__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14918__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14917__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14916__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14915__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14914__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14913__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14912__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14911__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14910__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14909__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14908__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14907__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14906__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14905__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14904__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14903__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14902__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14901__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14900__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14899__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14898__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14897__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14896__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14895__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14894__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14893__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14892__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14891__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14890__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14889__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14888__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14887__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14886__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14885__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14884__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14883__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14882__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14881__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14880__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14879__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14878__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14877__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14876__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14875__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14874__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14873__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14872__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14871__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14870__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14869__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14868__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14867__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14866__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14865__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14864__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14863__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14862__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14861__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14860__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14859__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14858__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14857__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14856__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14855__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14854__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14853__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14852__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14851__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14850__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14849__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14848__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14847__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14846__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14845__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14844__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14843__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14842__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14841__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14840__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14839__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14838__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14837__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14836__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14835__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14834__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14833__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14832__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14831__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14830__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14829__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14828__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14827__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14826__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14825__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14824__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14823__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14822__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14821__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14820__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14819__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14818__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14817__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14816__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14815__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14814__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14813__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14812__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14811__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14810__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14809__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14808__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14807__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14806__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14805__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14804__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14803__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14802__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14801__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14800__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14799__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14798__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14797__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14796__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14795__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14794__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14793__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14792__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14791__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14790__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14789__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14788__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14787__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14786__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14785__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14784__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14783__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14782__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14781__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14780__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14779__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14778__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14777__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14776__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14775__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14774__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14773__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14772__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14771__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14770__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14769__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14768__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14767__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14766__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14765__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14764__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14763__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14762__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14761__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14760__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14759__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14758__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14757__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14756__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14755__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14754__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14753__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14752__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14751__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14750__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14749__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14748__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14747__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14746__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14745__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14744__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14743__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14742__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14741__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14740__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14739__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14738__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14737__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14736__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14735__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14734__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14733__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14732__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14731__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14730__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14729__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14728__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14727__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14726__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14725__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14724__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14723__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14722__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14721__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14720__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14719__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14718__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14717__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14716__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14715__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14714__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14713__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14712__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14711__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14710__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14709__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14708__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14707__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14706__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14705__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14704__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14703__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14702__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14701__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14700__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14699__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14698__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14697__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14696__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14695__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14694__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14693__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14692__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14691__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14690__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14689__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14688__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14687__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14686__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14685__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14684__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14683__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14682__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14681__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14680__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14679__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14678__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14677__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14676__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14675__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14674__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14673__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14672__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14671__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14670__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14669__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14668__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14667__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14666__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14665__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14664__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14663__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14662__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14661__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14660__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14659__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14658__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14657__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14656__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14655__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14654__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14653__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14652__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14651__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14650__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14649__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14648__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14647__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14646__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14645__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14644__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14643__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14642__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14641__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14640__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14639__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14638__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14637__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14636__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14635__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14634__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14633__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14632__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14631__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14630__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14629__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14628__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14627__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14626__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14625__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14624__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14623__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14622__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14621__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14620__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14619__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14618__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14617__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14616__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14615__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14614__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14613__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14612__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14611__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14610__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14609__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14608__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14607__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14606__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14605__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14604__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14603__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14602__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14601__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14600__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14599__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14598__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14597__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14596__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14595__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14594__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14593__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14592__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14591__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14590__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14589__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14588__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14587__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14586__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14585__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14584__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14583__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14582__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14581__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14580__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14579__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14578__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14577__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14576__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14575__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14574__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14573__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14572__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14571__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14570__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14569__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14568__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14567__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14566__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14565__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14564__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14563__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14562__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14561__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14560__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14559__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14558__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14557__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14556__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14555__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14554__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14553__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14552__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14551__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14550__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14549__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14548__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14547__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14546__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14545__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14544__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14543__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14542__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14541__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14540__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14539__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14538__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14537__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14536__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14535__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14534__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14533__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14532__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14531__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14530__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14529__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14528__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14527__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14526__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14525__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14524__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14523__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14522__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14521__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14520__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14519__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14518__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14517__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14516__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14515__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14514__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14513__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14512__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14511__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14510__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14509__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14508__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14507__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14506__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14505__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14504__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14503__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14502__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14501__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14500__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14499__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14498__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14497__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14496__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14495__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14494__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14493__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14492__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14491__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14490__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14489__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14488__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14487__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14486__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14485__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14484__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14483__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14482__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14481__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14480__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14479__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14478__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14477__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14476__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14475__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14474__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14473__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14472__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14471__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14470__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14469__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14468__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14467__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14466__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14465__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14464__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14463__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14462__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14461__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14460__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14459__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14458__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14457__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14456__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14455__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14454__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14453__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14452__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14451__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14450__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14449__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14448__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14447__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14446__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14445__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14444__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14443__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14442__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14441__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14440__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14439__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14438__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14437__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14436__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14435__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14434__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14433__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14432__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14431__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14430__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14429__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14428__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14427__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14426__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14425__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14424__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14423__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14422__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14421__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14420__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14419__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14418__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14417__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14416__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14415__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14414__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14413__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14412__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14411__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14410__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14409__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14408__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14407__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14406__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14405__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14404__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14403__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14402__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14401__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14400__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14399__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14398__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14397__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14396__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14395__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14394__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14393__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14392__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14391__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14390__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14389__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14388__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14387__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14386__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14385__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14384__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14383__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14382__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14381__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14380__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14379__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14378__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14377__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14376__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14375__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14374__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14373__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14372__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14371__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14370__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14369__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14368__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14367__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14366__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14365__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14364__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14363__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14362__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14361__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14360__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14359__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14358__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14357__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14356__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14355__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14354__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14353__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14352__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14351__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14350__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14349__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14348__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14347__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14346__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14345__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14344__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14343__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14342__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14341__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14340__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14339__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14338__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14337__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14336__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14335__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14334__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14333__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14332__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14331__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14330__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14329__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14328__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14327__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14326__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14325__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14324__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14323__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14322__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14321__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14320__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14319__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14318__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14317__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14316__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14315__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14314__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14313__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14312__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14311__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14310__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14309__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14308__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14307__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14306__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14305__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14304__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14303__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14302__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14301__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14300__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14299__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14298__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14297__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14296__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14295__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14294__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14293__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14292__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14291__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14290__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14289__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14288__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14287__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14286__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14285__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14284__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14283__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14282__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14281__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14280__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14279__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14278__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14277__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14276__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14275__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14274__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14273__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14272__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14271__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14270__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14269__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14268__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14267__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14266__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14265__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14264__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14263__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14262__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14261__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14260__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14259__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14258__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14257__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14256__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14255__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14254__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14253__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14252__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14251__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14250__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14249__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14248__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14247__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14246__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14245__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14244__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14243__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14242__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14241__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14240__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14239__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14238__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14237__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14236__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14235__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14234__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14233__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14232__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14231__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14230__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14229__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14228__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14227__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14226__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14225__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14224__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14223__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14222__CLK (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15821__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15313__CLKN (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15312__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15311__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15310__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15309__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15308__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15307__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15306__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15305__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15304__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15303__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15302__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15301__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15300__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15299__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15298__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15297__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15296__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15295__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15294__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15293__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15292__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15291__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15290__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15289__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15288__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15287__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15286__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15285__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15284__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15283__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15282__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15281__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15280__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15279__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15278__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15277__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15276__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15275__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15274__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15273__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15272__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15271__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15270__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15269__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15268__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15267__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15266__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15265__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15264__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15263__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15262__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15261__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15260__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15259__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15258__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15257__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15256__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15255__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15254__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15253__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15252__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15251__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15250__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15249__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15248__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15247__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15246__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15245__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15244__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15243__CLK (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13425__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13422__B (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12835__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09097__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output6_I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_150_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_166_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_166_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_166_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_171_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_172_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_173_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_175_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_175_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_177_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_178_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_178_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_178_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_179_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_181_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_181_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_181_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_181_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_181_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_181_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_181_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_181_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_182_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_182_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_182_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_182_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_182_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_183_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_183_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_183_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_184_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_184_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_184_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_184_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_184_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_184_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_184_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_184_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_184_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_185_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_185_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_185_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_185_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_185_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_185_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_185_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_185_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_185_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_185_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_185_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_186_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_186_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_186_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_186_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_186_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_186_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_186_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_186_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_187_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_187_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_187_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_187_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_187_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_187_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_187_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_187_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_187_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_188_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_188_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_188_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_188_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_188_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_188_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_188_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_188_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_189_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_189_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_189_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_189_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_189_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_189_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_189_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_189_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_189_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_189_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_189_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_189_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_189_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_190_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_190_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_190_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_190_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_190_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_190_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_190_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_190_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_190_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_190_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_190_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_190_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_190_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_190_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_190_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_191_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_191_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_191_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_191_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_191_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_191_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_191_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_191_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_192_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_192_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_192_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_192_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_192_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_192_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_192_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_192_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_192_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_192_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_192_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_193_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_193_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_193_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_193_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_193_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_193_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_193_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_193_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_193_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_193_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_193_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_193_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_194_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_194_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_194_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_194_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_194_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_194_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_194_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_194_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_194_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_196_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_196_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_196_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_196_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_196_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_196_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_196_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_196_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_196_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_196_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_196_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_197_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_197_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_197_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_197_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_197_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_197_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_197_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_198_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_198_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_198_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_198_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_198_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_198_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_198_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_198_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_198_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_199_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_199_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_199_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_199_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_199_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_199_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_200_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_200_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_200_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_200_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_200_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_200_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_200_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_200_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_200_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_200_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_200_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_200_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_200_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_200_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_200_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_201_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_201_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_201_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_201_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_201_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_201_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_202_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_202_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_202_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_202_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_202_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_202_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_202_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_202_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_202_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_202_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_203_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_203_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_203_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_203_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_203_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_203_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_203_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_204_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_204_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_204_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_204_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_204_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_204_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_204_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_204_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_204_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_205_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_205_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_205_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_205_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_205_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_205_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_205_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_205_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_205_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_205_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_205_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_206_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_206_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_206_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_206_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_206_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_206_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_206_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_206_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_206_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_206_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_206_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_206_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_206_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_206_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_206_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_206_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_207_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_207_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_207_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_207_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_207_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_207_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_207_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_207_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_207_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_207_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_207_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_207_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_207_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_207_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_208_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_208_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_208_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_208_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_208_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_208_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_208_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_208_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_208_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_208_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_209_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_209_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_209_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_209_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_209_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_210_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_210_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_210_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_210_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_210_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_210_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_210_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_210_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_210_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_210_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_210_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_210_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_210_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_210_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_210_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_211_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_211_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_211_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_211_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_211_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_212_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_212_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_212_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_212_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_212_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_212_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_212_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_212_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_212_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_212_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_212_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_212_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_212_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_212_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_212_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_212_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_213_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_213_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_213_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_213_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_213_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_213_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_213_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_214_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_214_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_214_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_214_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_214_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_214_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_214_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_214_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_214_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_214_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_214_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_214_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_214_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_214_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_214_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_214_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_215_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_215_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_215_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_215_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_215_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_215_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_216_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_216_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_216_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_216_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_216_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_216_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_216_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_216_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_216_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_216_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_216_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_216_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_216_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_216_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_217_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_217_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_217_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_217_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_217_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_217_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_217_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_217_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_217_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_217_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_217_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_217_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_218_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_218_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_218_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_218_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_218_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_218_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_218_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_218_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_218_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_218_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_219_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_219_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_219_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_219_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_219_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_219_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_219_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_220_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_220_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_220_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_220_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_220_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_220_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_220_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_220_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_221_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_221_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_221_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_221_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_221_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_221_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_221_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_222_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_222_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_222_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_222_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_222_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_222_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_222_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_222_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_222_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_222_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_222_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_223_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_223_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_223_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_223_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_223_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_223_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_223_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_224_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_224_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_224_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_224_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_224_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_224_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_224_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_224_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_225_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_225_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_225_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_225_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_225_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_225_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_225_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_226_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_226_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_226_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_226_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_226_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_226_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_226_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_226_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_226_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_226_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_226_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_226_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_226_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_226_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_226_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_226_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_227_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_227_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_227_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_227_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_227_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_227_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_227_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_227_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_227_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_227_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_228_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_228_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_228_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_228_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_228_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_228_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_228_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_228_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_228_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_228_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_228_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_228_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_228_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_228_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_228_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_228_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_228_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_228_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_229_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_229_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_229_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_230_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_230_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_230_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_230_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_230_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_230_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_230_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_230_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_231_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_231_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_231_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_231_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_231_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_231_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_231_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_231_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_231_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_231_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_231_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_232_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_232_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_232_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_232_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_232_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_232_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_232_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_232_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_232_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_232_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_232_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_232_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_232_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_232_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_233_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_233_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_233_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_233_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_233_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_233_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_233_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_233_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_233_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_233_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_233_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_234_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_234_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_234_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_234_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_234_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_234_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_234_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_234_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_234_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_235_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_235_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_235_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_235_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_235_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_235_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_235_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_235_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_236_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_236_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_236_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_236_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_236_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_236_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_236_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_236_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_236_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_237_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_237_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_237_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_237_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_238_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_238_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_238_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_238_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_238_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_238_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_239_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_239_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_239_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_239_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_239_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_239_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_239_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_240_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_240_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_240_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_241_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_242_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_242_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_242_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_242_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_243_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_244_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_244_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_244_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_247_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_247_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_248_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_248_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_248_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_248_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_249_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_249_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_250_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_250_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_250_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_250_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_251_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_251_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_252_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_252_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_252_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_252_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_253_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_253_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_254_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_254_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_254_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_254_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_255_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_255_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_256_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_256_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_256_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_256_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_257_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_257_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_258_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_258_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_258_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_258_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_259_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_259_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_260_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_260_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_260_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_260_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_261_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_261_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_262_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_262_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_262_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_262_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_263_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_263_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_264_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_264_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_264_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_264_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_265_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_265_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_266_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_266_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_266_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_266_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_266_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_266_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_266_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_266_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_266_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_266_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_266_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_266_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_266_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_266_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_266_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_266_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_266_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_266_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_266_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_266_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_266_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_266_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_266_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_266_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_266_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_266_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_266_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_266_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_266_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_266_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_1365 ();
 assign io_oeb[0] = net8;
 assign io_oeb[10] = net18;
 assign io_oeb[11] = net19;
 assign io_oeb[12] = net20;
 assign io_oeb[13] = net21;
 assign io_oeb[14] = net22;
 assign io_oeb[15] = net23;
 assign io_oeb[16] = net24;
 assign io_oeb[17] = net25;
 assign io_oeb[18] = net26;
 assign io_oeb[19] = net27;
 assign io_oeb[1] = net9;
 assign io_oeb[20] = net28;
 assign io_oeb[21] = net29;
 assign io_oeb[22] = net30;
 assign io_oeb[23] = net31;
 assign io_oeb[24] = net32;
 assign io_oeb[25] = net33;
 assign io_oeb[26] = net34;
 assign io_oeb[27] = net35;
 assign io_oeb[28] = net36;
 assign io_oeb[29] = net37;
 assign io_oeb[2] = net10;
 assign io_oeb[30] = net38;
 assign io_oeb[31] = net39;
 assign io_oeb[32] = net40;
 assign io_oeb[33] = net41;
 assign io_oeb[34] = net42;
 assign io_oeb[35] = net43;
 assign io_oeb[36] = net44;
 assign io_oeb[37] = net45;
 assign io_oeb[3] = net11;
 assign io_oeb[4] = net12;
 assign io_oeb[5] = net13;
 assign io_oeb[6] = net14;
 assign io_oeb[7] = net15;
 assign io_oeb[8] = net16;
 assign io_oeb[9] = net17;
 assign io_out[0] = net46;
 assign io_out[10] = net56;
 assign io_out[11] = net57;
 assign io_out[12] = net58;
 assign io_out[15] = net59;
 assign io_out[16] = net60;
 assign io_out[17] = net61;
 assign io_out[18] = net62;
 assign io_out[19] = net63;
 assign io_out[1] = net47;
 assign io_out[20] = net64;
 assign io_out[21] = net65;
 assign io_out[22] = net66;
 assign io_out[23] = net67;
 assign io_out[24] = net68;
 assign io_out[25] = net69;
 assign io_out[26] = net70;
 assign io_out[27] = net71;
 assign io_out[28] = net72;
 assign io_out[29] = net73;
 assign io_out[2] = net48;
 assign io_out[30] = net74;
 assign io_out[31] = net75;
 assign io_out[32] = net76;
 assign io_out[33] = net77;
 assign io_out[34] = net78;
 assign io_out[35] = net79;
 assign io_out[36] = net80;
 assign io_out[37] = net81;
 assign io_out[3] = net49;
 assign io_out[4] = net50;
 assign io_out[5] = net51;
 assign io_out[6] = net52;
 assign io_out[7] = net53;
 assign io_out[8] = net54;
 assign io_out[9] = net55;
 assign la_data_out[0] = net82;
 assign la_data_out[10] = net92;
 assign la_data_out[11] = net93;
 assign la_data_out[12] = net94;
 assign la_data_out[13] = net95;
 assign la_data_out[14] = net96;
 assign la_data_out[15] = net97;
 assign la_data_out[16] = net98;
 assign la_data_out[17] = net99;
 assign la_data_out[18] = net100;
 assign la_data_out[19] = net101;
 assign la_data_out[1] = net83;
 assign la_data_out[20] = net102;
 assign la_data_out[21] = net103;
 assign la_data_out[22] = net104;
 assign la_data_out[23] = net105;
 assign la_data_out[24] = net106;
 assign la_data_out[25] = net107;
 assign la_data_out[26] = net108;
 assign la_data_out[27] = net109;
 assign la_data_out[28] = net110;
 assign la_data_out[29] = net111;
 assign la_data_out[2] = net84;
 assign la_data_out[30] = net112;
 assign la_data_out[31] = net113;
 assign la_data_out[32] = net114;
 assign la_data_out[33] = net115;
 assign la_data_out[34] = net116;
 assign la_data_out[35] = net117;
 assign la_data_out[36] = net118;
 assign la_data_out[37] = net119;
 assign la_data_out[38] = net120;
 assign la_data_out[39] = net121;
 assign la_data_out[3] = net85;
 assign la_data_out[40] = net122;
 assign la_data_out[41] = net123;
 assign la_data_out[42] = net124;
 assign la_data_out[43] = net125;
 assign la_data_out[44] = net126;
 assign la_data_out[45] = net127;
 assign la_data_out[46] = net128;
 assign la_data_out[47] = net129;
 assign la_data_out[48] = net130;
 assign la_data_out[49] = net131;
 assign la_data_out[4] = net86;
 assign la_data_out[50] = net132;
 assign la_data_out[51] = net133;
 assign la_data_out[52] = net134;
 assign la_data_out[53] = net135;
 assign la_data_out[54] = net136;
 assign la_data_out[55] = net137;
 assign la_data_out[56] = net138;
 assign la_data_out[57] = net139;
 assign la_data_out[58] = net140;
 assign la_data_out[59] = net141;
 assign la_data_out[5] = net87;
 assign la_data_out[60] = net142;
 assign la_data_out[61] = net143;
 assign la_data_out[62] = net144;
 assign la_data_out[63] = net145;
 assign la_data_out[6] = net88;
 assign la_data_out[7] = net89;
 assign la_data_out[8] = net90;
 assign la_data_out[9] = net91;
 assign user_irq[0] = net146;
 assign user_irq[1] = net147;
 assign user_irq[2] = net148;
 assign wbs_ack_o = net149;
 assign wbs_dat_o[0] = net150;
 assign wbs_dat_o[10] = net160;
 assign wbs_dat_o[11] = net161;
 assign wbs_dat_o[12] = net162;
 assign wbs_dat_o[13] = net163;
 assign wbs_dat_o[14] = net164;
 assign wbs_dat_o[15] = net165;
 assign wbs_dat_o[16] = net166;
 assign wbs_dat_o[17] = net167;
 assign wbs_dat_o[18] = net168;
 assign wbs_dat_o[19] = net169;
 assign wbs_dat_o[1] = net151;
 assign wbs_dat_o[20] = net170;
 assign wbs_dat_o[21] = net171;
 assign wbs_dat_o[22] = net172;
 assign wbs_dat_o[23] = net173;
 assign wbs_dat_o[24] = net174;
 assign wbs_dat_o[25] = net175;
 assign wbs_dat_o[26] = net176;
 assign wbs_dat_o[27] = net177;
 assign wbs_dat_o[28] = net178;
 assign wbs_dat_o[29] = net179;
 assign wbs_dat_o[2] = net152;
 assign wbs_dat_o[30] = net180;
 assign wbs_dat_o[31] = net181;
 assign wbs_dat_o[3] = net153;
 assign wbs_dat_o[4] = net154;
 assign wbs_dat_o[5] = net155;
 assign wbs_dat_o[6] = net156;
 assign wbs_dat_o[7] = net157;
 assign wbs_dat_o[8] = net158;
 assign wbs_dat_o[9] = net159;
endmodule

