magic
tech gf180mcuC
magscale 1 5
timestamp 1670237842
<< obsm1 >>
rect 672 1538 69328 58438
<< obsm2 >>
rect 2238 345 69874 58427
<< metal3 >>
rect 69800 57792 70000 57848
rect 69800 53816 70000 53872
rect 69800 49840 70000 49896
rect 69800 45864 70000 45920
rect 69800 41888 70000 41944
rect 69800 37912 70000 37968
rect 69800 33936 70000 33992
rect 69800 29960 70000 30016
rect 69800 25984 70000 26040
rect 69800 22008 70000 22064
rect 69800 18032 70000 18088
rect 69800 14056 70000 14112
rect 69800 10080 70000 10136
rect 69800 6104 70000 6160
rect 69800 2128 70000 2184
<< obsm3 >>
rect 2233 57878 69879 58422
rect 2233 57762 69770 57878
rect 2233 53902 69879 57762
rect 2233 53786 69770 53902
rect 2233 49926 69879 53786
rect 2233 49810 69770 49926
rect 2233 45950 69879 49810
rect 2233 45834 69770 45950
rect 2233 41974 69879 45834
rect 2233 41858 69770 41974
rect 2233 37998 69879 41858
rect 2233 37882 69770 37998
rect 2233 34022 69879 37882
rect 2233 33906 69770 34022
rect 2233 30046 69879 33906
rect 2233 29930 69770 30046
rect 2233 26070 69879 29930
rect 2233 25954 69770 26070
rect 2233 22094 69879 25954
rect 2233 21978 69770 22094
rect 2233 18118 69879 21978
rect 2233 18002 69770 18118
rect 2233 14142 69879 18002
rect 2233 14026 69770 14142
rect 2233 10166 69879 14026
rect 2233 10050 69770 10166
rect 2233 6190 69879 10050
rect 2233 6074 69770 6190
rect 2233 2214 69879 6074
rect 2233 2098 69770 2214
rect 2233 350 69879 2098
<< metal4 >>
rect 2224 1538 2384 58438
rect 4474 1538 4634 58438
rect 6724 1538 6884 58438
rect 8974 1538 9134 58438
rect 11224 1538 11384 58438
rect 13474 1538 13634 58438
rect 15724 1538 15884 58438
rect 17974 1538 18134 58438
rect 20224 1538 20384 58438
rect 22474 1538 22634 58438
rect 24724 1538 24884 58438
rect 26974 1538 27134 58438
rect 29224 1538 29384 58438
rect 31474 1538 31634 58438
rect 33724 1538 33884 58438
rect 35974 1538 36134 58438
rect 38224 1538 38384 58438
rect 40474 1538 40634 58438
rect 42724 1538 42884 58438
rect 44974 1538 45134 58438
rect 47224 1538 47384 58438
rect 49474 1538 49634 58438
rect 51724 1538 51884 58438
rect 53974 1538 54134 58438
rect 56224 1538 56384 58438
rect 58474 1538 58634 58438
rect 60724 1538 60884 58438
rect 62974 1538 63134 58438
rect 65224 1538 65384 58438
rect 67474 1538 67634 58438
<< obsm4 >>
rect 42966 1508 44944 49607
rect 45164 1508 47194 49607
rect 47414 1508 49444 49607
rect 49664 1508 51694 49607
rect 51914 1508 53944 49607
rect 54164 1508 56194 49607
rect 56414 1508 58444 49607
rect 58664 1508 60694 49607
rect 60914 1508 62944 49607
rect 63164 1508 65194 49607
rect 65414 1508 67444 49607
rect 67664 1508 68866 49607
rect 42966 345 68866 1508
<< labels >>
rlabel metal3 s 69800 2128 70000 2184 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 69800 6104 70000 6160 6 io_in[1]
port 2 nsew signal input
rlabel metal3 s 69800 10080 70000 10136 6 io_in[2]
port 3 nsew signal input
rlabel metal3 s 69800 14056 70000 14112 6 io_in[3]
port 4 nsew signal input
rlabel metal3 s 69800 18032 70000 18088 6 io_in[4]
port 5 nsew signal input
rlabel metal3 s 69800 41888 70000 41944 6 io_oeb[0]
port 6 nsew signal output
rlabel metal3 s 69800 45864 70000 45920 6 io_oeb[1]
port 7 nsew signal output
rlabel metal3 s 69800 49840 70000 49896 6 io_oeb[2]
port 8 nsew signal output
rlabel metal3 s 69800 53816 70000 53872 6 io_oeb[3]
port 9 nsew signal output
rlabel metal3 s 69800 57792 70000 57848 6 io_oeb[4]
port 10 nsew signal output
rlabel metal3 s 69800 22008 70000 22064 6 io_out[0]
port 11 nsew signal output
rlabel metal3 s 69800 25984 70000 26040 6 io_out[1]
port 12 nsew signal output
rlabel metal3 s 69800 29960 70000 30016 6 io_out[2]
port 13 nsew signal output
rlabel metal3 s 69800 33936 70000 33992 6 io_out[3]
port 14 nsew signal output
rlabel metal3 s 69800 37912 70000 37968 6 io_out[4]
port 15 nsew signal output
rlabel metal4 s 2224 1538 2384 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 6724 1538 6884 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 11224 1538 11384 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 15724 1538 15884 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 20224 1538 20384 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 24724 1538 24884 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 29224 1538 29384 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 33724 1538 33884 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 38224 1538 38384 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 42724 1538 42884 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 47224 1538 47384 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 51724 1538 51884 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 56224 1538 56384 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 60724 1538 60884 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 65224 1538 65384 58438 6 vdd
port 16 nsew power bidirectional
rlabel metal4 s 4474 1538 4634 58438 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 8974 1538 9134 58438 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 13474 1538 13634 58438 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 17974 1538 18134 58438 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 22474 1538 22634 58438 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 26974 1538 27134 58438 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 31474 1538 31634 58438 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 35974 1538 36134 58438 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 40474 1538 40634 58438 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 44974 1538 45134 58438 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 49474 1538 49634 58438 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 53974 1538 54134 58438 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 58474 1538 58634 58438 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 62974 1538 63134 58438 6 vss
port 17 nsew ground bidirectional
rlabel metal4 s 67474 1538 67634 58438 6 vss
port 17 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 70000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 28066146
string GDS_FILE /home/runner/work/gf180-mpw0-serv/gf180-mpw0-serv/openlane/serv_0/runs/22_12_05_10_54/results/signoff/serv_0.magic.gds
string GDS_START 22272362
<< end >>

